PK   ���X��/�   ί    cirkitFile.json�]m��6��+��`y�����d7� ���r��0�%�����u�3��߯(�m[�l�����f�gZ䣇�b��"��N��O�z��l��O��i�YO�J;�|(�է���b:y\����o�����������:Yl�Zl��<��Z�V%��DbLV$y!ʤ4�ɚ��������}���~�Fs���Es���Es���Es���Es���E�́� �!��?n>��d[�bd���C�]�~I���&��d����Yn>>n��z7�e���")��ILS.�ҖYR)-�]�&M���L�9���o����L}��P��'f�$`� ���C��6���lb��?�Ă?��!�aC��|b�5��A,�FT�!�����lb���lb���S�mg��\��M�¹�n�����mzq��s[��Z��[Pp[��K��u�.Q��ă:�ļ��܈��I,;�eG� Vv+;(;�eGڏ�����Nbى���Ncee'����`eg�����Xvbn���X�A�I,;1O��K�����Xv�|!�+;(;o���[�� OT9V�9V�Pv�g��j��eS�D�K���I�P�lѨ��u�ьZ0�^`�^`�[PR�%�-�
$ħ��1����@ď���!:�UUIpX��'���9�Za�I0?��,?px��'���gG���!���sL���YX~��}��ja�I0?��,?p���'����u�������s������O���-`���,?	��6c��������?�[8�x�y��;^pt ��/��+l���s�S\��G��,?	�����~��$��ۜ�8���`~n[X~���O���a`���,?y���������w7"�ɫ��=<�zw�����}��w7�����9�zw�����CՆ�vL������<����L�����>�H���L��q�ϵ{L��z��H(������v��{���g��Y�kOSp^_p_�r^��#O���EeKc�H��^$��:ɕ�2V-�F�iQ\�w��3��?죪��:E#�y�R,#I�ԉ�7[�(�!E��m��������m���l{��U���K�3k�DɬN��uR�N��X.�ʦ�}��P��^Y�x�z�dm3=�^�Y��MA������T��*K��0��h�y3�Ѻ��Q���X��y�UO�#���f�y�伹`GU��Q��}�ȡ[�Qa��������F�Y�r%t���?��n����&q�0�Ε(4�>s�\�B��3��(4�\3g]0U��˱�̦�4�Qi��˸�̡d�C�0��a%�J�9�l߄b*��e^%�Q��{�&e��DS�UW��Z6����y�Q���"y3�\���HޜWS�?��v����͖�Mq�h�L��IP��c���� ��FF �6��0�
���y0�@@m5�B�ŗ_��(��M��1�Q�
�T��hx�
��lm�7� L$�j��6�nK��F!�X'��0�Bڇ� N0�-a���A�`6\�l��!�@�`v\��o�>�"����9�0;�`v|�ğ��)A��1�'Aq: �uV39���)-s����}�B'�W0;�B�'1q�A�4����U�~�C8*�����
��\��	t��Q�r���#��a58*P�cp�s'b$�=�G�u�~^E�����@����Ϲ��@��(�1���1�G���:W?Wc(F�']�ȵ{X#�1���1r�_�ȵ{�#���"�ϖ���	��� �g��(l�Hَv�wy��Hَz��6�I���8��(lY�Hَ���6�����8a�(l��Hَ���6�����8��(lY�Hَ���6�����li A_ Ɖ˼���o �|
�m S$)�q�Q��H�a����8q��������V3
�@�H<,R���e���[/�"H���e��$�	a���K��8q�(l9%�Hَ���6�o���8q�(l�(�Hَ�E����ҳ�{x�J J����9,(=���g��������ҳ���l�����#&��}���ȋ����p߱�;�e"�F����ܑAs���A�;2b�N�ޑ��(�����#ߥ��x�#oe���'��M-��F	@�p�9�bST^G��T	@�)�ؼ� �\nN���,o�D洜|�4��ֱ�)i�	�Ħ�t\j+��b��2=-�My]��� (�\b�;�rSwc�5PnN�������L� .7}�輌ׇct�E���7:�b���l0|;R�N����(��H%:�" F�0w�F�1�1e0c���g��&"`0c�`Ɣ��)�S3��A��ja90��|�E&6��u2�9_���>��]HG���w����}�@{���M!�@@{?����!�@@{�����!�@@�� ���1 �@@�x�t�}0&g�qff�%�p��!��vK��F!�O'���0�B:��N0.aF�t�1�`v\��8
鐎�	��p�W0;�B:�#�p��q��(�C:B'�W0;�B:�#�p��q��}H�t�h���D j !�5���
��\�!��3�Q�r�k !D�Y&4*P�cp�#�H�;ǄF�u��t�	xg�Ш@���5��"��(�1��B$��]B��:�@:B��sKhT�\��HG��wf	�
��\�1�8����Ïr��6�����Ha�8q������8��(lC��Hَ~��6�����8!�(lC��Hَ���6�����8��(lC��Hَ���6�����8!�(lC��Hَ���6�����0N\6
�P:B8,R���e���#��"e;�'�q�2?�)�q�Q؆��a��'.�m(!)�q�Q؆��a��'.�m(!)�q�Q؆��a��'.�m(!)�q�(�w�#����#!�g����(={��HG�G���{G:B>J���{�`0��w�t� �����'! ��}ǆ�IG�z-�;OsO:B F���ܓ� �����#�`�Xc�X����t�|��*:�U��t�|��r�NG�G��妙�NGx%6!�fE�#���������rSw���Qn�nt:B>��	2:!������u ��h��H%>! ���#��t� �ߎT���F�5����1�1e0cʀ�̘2�1e0c�`Ɣ��)��b��b{S����Qι|��_&Gq���W�ϓ��N'�V��i��P.�j�Z�7۪�N޾{�p29��?N�3�Ϋ{�}���H��Ͳ��\�,ыE��/����$�)Im��*S�6�0Ἒ�w��ՑQ!ǟ�ys���	C{^iH���HK8FWǮȝ����3��+�k]��zs�V��o�y�ޜ�F�q���6�Yv����a4!��YT:����uŮ�U�K�)��fK氾����t�t�#=n<����љ��7?�7_���c��8R�������������?��~�f�[|�E����1��������g���O���Ѯ�XZ��w���,��p��2x����^eE�$�N\����7���,���:^m�4��7X1��/�BHp�O��	��`�ϵ��o�~y����Q��������ˈ^�ưB/NCL'|��
�T�o�^g���!�q:�x^�_n�|���i���
��U��s�s���]�Ll���m&6�~�7�b�k�ɂ��u�d����Zg�`C�w���?��He|R�GJ0C��O��I�<R��	����!,/��l�_>������J��c�Mpy l�a>������J��� ���.�yU G��q� ����"�Y�=U {�bt�Nͤ0�-F��b�X����dLZ ��bth�LZ [��8\t����
`�}��Y��̸8�}Z+^�K�_��JD~X~�k*���2��� ���\G�l������_��If{�L�8<�����K2��e���A���F��^/�,"?,��u���zYeqx�a������<��^"Y�8����c�n�숓�7p-$S�^�Xf�=~��K<��FG+�͊\��cx�3#Rx �`�!:��Obd�c�C�:12D�2`�������0��%�@@��!�a�2F  F���0t�"#Cthf�\��!:�3]����0te"wM��rW�џY�C�"12D�)`������?�����@  F��k�1x������@�H�a����ޔ;$��b���@G1`�������0���@@��Q�a�*B  F��(�0t� #Cts������nۡ9_���ݭC�"b�������X���9���sr`}o�����Nš��V@��V�pu�?"2������᩟� \E��/�D\M�O�jb`��`��~�o(WO�=�C�z��-{Ҟ���wmG��������G_�ǩ�}��A}�_O����8���?��>N}n��Lf���Տ���3�z�F��ׁ�I#}Y_�'QE��}8N¯+�}q����N��}@�\�����8��L~�W�ō���8t�8l��������X�������:����k�E�}}, ��^,�o�cp��Z`_G-Xv�K�pG��s�K��|���;4wh��0ܡa&\s���
�E_�G/��=�������\F1�r)�b���wg�<����Y�̈́.�t�����:@k5����~0n7���K�+��𖮂t5���ZlW����&ls�*WC���h�jWC�{�&1�O�*��	��v ��	�*�8�b�����oi�ߌ�k\]Ӿ��5��qu����5��u5���&1�{�r��罒����9=$��ZKW���A�dL�W����P�d^�?���ټ���me�a_�/Åټ����B���6��(g1�"�/w��/�u�x�_��G�k��Y��,��w�e{��;&C��{��Dހ�_��l�1D���/2|f⓻�st?����y]�.��K�{���yd����Y��:<R�#}x��G��Q�?��2�Q~x����ã�{�.��M��q��ǖI�i��4�M�(}Aʣ e@�G��z����L�W�f3X=휆�Z+]�:Y�:O�"͓�
�Ժ��,���y��j����z�H]̊�?�m�|~t�E��kq�J=(iZ,������ed<��ܹH���W�o7��v���p�����pC����ۮ��΁u����=�N~*�ݿ~��_im�4�y�"���Ӈͧ��_��mS><�����u��Z<�/����x^m�j�vGԩ�>��g��w�[wOf?��bg\��߿y^�2���jC�x����hD���E�٩�����S�WN����-ALd�K�U2�K΋\f��dI6'+t�뺞���_��S�*9���O�r��E����f�"�rOw�P7;���.�C?SD63gj�����i��*��Y
v��KZa�B�g�Tevv�����S�:$Rk]�w"�����s�ڼ�z"gz�i�r�1k-�o��_Ve�}^��|���]jZ%��f)Ţ���,��u�\�.DSWIaK���`��e�\�n�f��"J�z�z���K-4J�g�,��gbfi�����%_:}M�M��s �m�YfOs���L]�q�'=�	qAVF'n�'��]	�H����f�]�'Q+�]=�6�֞����(d�� ���eK���M���)/{����̨S�W=X,�C3��Ҵ������Nw��ɢc�UO�\ŕK�����3�4OXi.ʵB���p)q	f�`4S_�=�2�ջ`1�v�5X�ȘR*
K�`�"���`)�U�`)_u��|��(���b]��A��m_�4���+g��U�f�P����[�~�������n���d�~���߈TVº��ZT�IK}62�Z,�12Km���ǇM������n]2��&�,	@�$�/��$ot�TU�\�u[׽����_J��W^��)s�,��I�,e%�<K�޷����YeeK���&э#L�\����Ei�f�d�)�|�v�_���3���qV:������Yd�*��-(�W�ZRP�U*U֫Q|]n���w���%����&ɔ���)�.��,�����|��y��ٔ�h2%�D(��X�p�Z&J-HjbI̲C;���c��jW�M�����D_�P�,�{��/ߖ?m�>�7m��9j����7�ݗU�����>O��(;mVu@�f��Q�jr5�nKQ�[VK�ً��0�e�.��S�4-�e�l�bQ��BIR�&/���)�(\�}k�� �%͐�$�2�:���B�J6���*�]�Le�I�����IN���)51W�l�+�r�����6���S�{~�������7o���7��7�l���'o\�7�m=}�ۼ�>��l�UyK����-��f��X���m�X���z��l�����^�Z�iY���do=��-,}��ɩ���w���<�I��>��S��,��!P;w+i4�hҮD�d�Z�Di[�J��62.l���6$���0�/U��ӕy�Dz�唄;Ӆ���м����B��Ō����F�TR�K�*��u��OIs��N��FN�ϡ	��>R��9%�JmE�`v��s�t[���I�jQ���%�vQK�d��	u��lYg&[F)}������B�s�{����ȎkN|��\T-���*�3I�uq��E�H����L��ybt)h�!aE��"K���-mE��
��jݒU�3C�f���̸E�¾,0��!�	K�ס����� �T��vF�QV� ʤ3�'e�
���e�)�vh���Ϭ�RvfRuZ2�:?<Z�c1��אּ��¦\�`�G�rq���bd��V��b|zg&	-3G���)1��l�K1�QKQ�v��Pk�T��(	�L�0ϭ<k�3�B���h0�ff�Mi�>V3k��G�S����ܽ}�@�ȥ=p+���!M�O�dӅN��NŨQ2ϤJ��%S�j������Z����t��&�ұ�\��w�ŭ��p|�R�в]�$�E�Vl2��BѤabsM̌�X���u�q�R�؊�tmF��N�j�*ϲ�X��f۔8���:���@��-��i�R�Xh��F���V����k��Z���t��L��^l;Z�I��F�S�� �K��HM^u���RE)��H�mN��8.��r.�%�CzKRo��2����h���NO��#}l��Ѡ�N�#�&�D��b��HI�2yRZ���+�-��Ua,)}Nl~��s74�i$jb��v�mtYP��Z2�dwl�ٓr��$�[�LK�4��yh�����/b�w+'�����>,��#��HًSq{�w7��Փ݆�9IHg����OC�+�n�i?}ZU����L~��^��î��i�$�v��V����-��꫗O��o����O�C���g��b8
F� �ɰ��Ix��~�>��w�j����*T�&�j[~�I����c��Y�wߗ�-ů�'���w������|r�}����u$_Tm������
L��r{G)���R��Vd��7f�~��~�T��>���H��ۇ�S�,^}PC�Ov�����N]N�C�i/#���{��.��@��b�O�� C�C
�fH�f�1U���ew���R�P�R�.b�@��jPK��T���8հ2^5pC�Ɓ�@�h��Sw^�5/���-t�/J�<�R}6#���������.��U�(tqG�SvQ�2X�
�FZ�*]^U�{�D�G�9�[�q�<=/�����:VY���,ɥ����j �{J�n�>Q�7��{N� � Ql�d2��P5��܇�@wK���ᥔ�m0�T��,U�,���y�3���{���ܥ*��]8�j�t�S,U�bn�~p�x˒7v���,z<e��vEߧ,�DϢG�X���}X�K�*�̋/��n#�]Q�y�x�u�^m���<�_h槯3�-UG��J�=�+ta����9Ps��j��YE������`�9��9?��yM'�K����2w��{΍Bu�s�tDO�ܚ�0䙞�7�G�a8�9���=�x0�_���������_�պ�e���������"�������\5a��z�W3��/P���^����������N���/�|۔����wZ�.~3.��jY��H����b��K_��R�9�r�cl��V��R}�����w͟�]�]��2Ҩ������?�������ow�Gw��ݏN�������?�O����of���PK   ���XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   ���X� ���� 
� /   images/38cb4f51-bc72-4d24-b782-e5d855ce8001.png�|gX[n�c��"D���  M����t)���!�H�.���*��@@�tB(�	�����{�ϛ�<<g�^�]k�k���*�2�etMQAV�R	���"�˅�_������>��B Ǘ�*@@ �o�/Q���&�#���sGM�׎�/�MA���|�6�&/ߚ��ڛŭIЁ@�@���\�W&\]L��{Tw��_����(���i�m���?t]l���c���c}y0�"r��n>�~�2�4�܇���y���:]=�*���u:�����,V�;S8ܘ��`��������Q�x�_���YL�F���N�I���[̪��9���?-�%O�I��;�rv(Y�J�ӣ��7ǉN9.]^;sn���g��/~���7��w�矤��2�Oߒ�~f�s���&�`O�V��2������[�
�β�G�~�z,�x�T\�Bgv=�@�(��5������ЅM�9���<�T)V��m���q�X�
k����8k~Y�֖���Q=�AٗmYo� "�~A!�����K���WS���>�7��eO�r�D�ơW!ԁ����F�{�v�ٺI��G��h0ՙ]8jY����o�/8�\����q*���⩛6�萕t��嶋�Q��E����Ma��?|)�?�晬BuGQ¡S�wf0�'����򇞨�����?�����}oy�{x*��h����,���B�4�*���caH���%u<�@�a��%���{��PZ|g�$Ӑv��+�>F
Z|�[\�U��5���:��Gac���|�{I�5�݁(������Y"��S�ʨ)^Q/��β��抖��h��/�Jq�U�_��:\�K��I��\�pk�*	(���t��Rj_k��i�z8-o6"���<7��f$Rv?��&hD�K�ean��AO������5[�U�tB��&�lb5�53$f��K_�S�j�nl�C[A ���>��fQ��b9���	Ysl��^�䟧E	���"]`i�ePybГ�O��ݛqo���XZ�GXP��؂�J_�]�Mq&(O���������O��oW��4����L���T$mW̄��-�-��w�
S���<��f��p��)k���N�j)����s��y&D Z��!��5�G�D#=�g��B�*�kb�^m{b�R����P�xs�s=����� ���R^�j��)���h+�ݰ����oF��3q���#��W�Ev?��b#�Ќ�C^�,�U�4����2��A<�z!�P"Aѓ]���~#)Pz�:q���Z�z����A��Un���@W4������AK�WI��=�5���r@�+J�:e/_��&iК@om��*�2h��w�0*��;7(�#"p��{�갥LƇ����	ý�b����W���ވ��DA�?)^�k�d�\X0��;0�FM2�%/�u���go���ܖ�Yo�� BH B$�2E��o;���v�_9z�To��yK�b�mFrv����f��J ̴(CN�w-�)�zܞ�1�i�Z�3�i����Jl�Y�@,�Q�=�kI9�N:[�9Y�CznE=��ܓk�k]��l�q]G<�����T�D�P��@�[�I�қ̺��e|�������k����dr��r@�B��S�VIr%Պ:���B`�(�i���W�t@x�Dp�o�) ��jN���j���#��A�qN�U�8�cE�n68�S���3b�A�
;yTr�}�Ȏp�W�H,�j�b�#g3��)��`F/��qYh��i�/sD�/��kF)�h�4gy]h8�����q�Y��Mh&�$/)�j�7K�zpb�;˥�6��Q;���S�1�G<�?���ϣ I�I�4��t7����bn��:�q����6nDrvn�8�LVW=�0i�i�~��|�n'W�x<*�L�-2	6�eDZ�k���
c�@2�sŧ���#	.�X��c�X�;J����t�df�� �OS�U+��'�f��N�atn�ɒ�o"���
��Ū�A���"q�O�7z���5�:V}�>̐0�RB�@�
g����ӊ`2�9����L�fk@�R�wђ��B�z�_�04n";،K�N~�g��M-����?�?��8�Zo��U�~o��*yȩ�ʪ�#!���$���|I0f�g��
��[��W��s��t��a�rє��p��ӂ���a���z��ꅖ=��'`%�������^��2�	Z�)XKS��DS��U���LF��A��S�å�X�W�3����H���_�\�+x6�xN�3n&؃Z����Nշ08O|g�����L֪J����/~[0Th�r��T[���1�1�)?򥨧�D�RA��S�o
_�!Lv,���zk�21 ���~J_"�&�f�=S���Sw'�^�}�����lbm�ec	��=/�גU��T&�BK���+�t7���l��W��͡���D���,c
&]�=-����xUV̒� ��K�ˑ&0Wn��Ǖ��s ���*��� �f�I�$/�+p�{�T%�U��O]�&�d���i�\�yꉭ�9�-��"Zg	�*��dU-���Eh��oe'v�N
_��}d��g]0��c.~�R���H4_?�1sD����\EA'䢬�d�X=9�� g|�|��FDt�Q���6�B.ҥ:�w����ZZETyVͬ8��;:�s	0��hЋ����x��Q����8IR��<�Vv{t��Y?$�f���<�/
7���V���!D ��S�~�J�g[^����e/77 ����~�9��-�p��%!D	ܥ� �	FaYAwo��-��J1D6�	v�C�Ӓ�~�GP�(�m����W��m�rsr�S7#�MF��������yyy�ɋ�FjM��FK9˭�M��w'-SL�7B��_�/�.�<#��eRHG�8�(;� *h�B|��5g?���(�3�ȇ�'�;�8�>k0K
�L��1zI0���،��D�S�,O=F�;����T��-�9Z��n�]St�#�AB2��'��)ν����(S%��T���3M��k�U݋�5b�~VT�����4��e<4*%�\�㟣&,t��ds�ψ�]-�V0�r�����o�� �����SIb��Z�w��d������e�oie��bA���G̴�7>�=m_1�Y�yN�x����C٫��߿B����&�gP�<x4�
��OIIi��4�Xwk��u �<�W�_����C�-s��L�����xݣ�J>ս;��Vxhhcס7��v�N��������Q��L�ɿ"��٠$3'gGp��V��F�&Nl�-i��2,x�|w?i�6��v&D��S�O!hm���$�/|N=ӗف�ޤ$3�88 !\R'�j̀�K �L�">Q+�ZZN����1c3t��\}�������oIf�ۚeeeFIǎ�^;C�����!Bx���|Uz��P!�������%�*�ԙl����_���b�Ť?������1K1��f�f"����]�8�{�$��YW�K�aM$����C:�i�%!Ġ����n����ү]hi�Bլ�uBe)����w�rg��A����k��nP���ve�4w�.0WCU:cZ8����S�������inW�7���u����R�ʢRPd"'�;������ѯn��,�~�`Lf*����Ò7���
�n�l\`�GG���x��7=T��'�W�睘�S�q�B�ʥ�4�_^�5�E7����Y���0}�;r�C/v?�cY�5ag\��a��R(-T�4�������I���[k~�ͮ�<����a��I��Qx�����W!Vf>�{�mk����VlX���f��iz�K��x�x�ʣ;*��x2�t�����OK�� �뮥���N~d6	S<P>>;�3��!i��gj�5`�L�8��p���/:$!y�Fx��U�
�V�T�ZUB��F�w]�^�9��D� �OAqf�`����kג�����XN���f�Su��wW������N�� �#���z�wR�s�f���KC�ڿ��M3���z*���e�I"B�	"B�f�,�Sb�,�jsxHa���rJ����ؼ�^Kq�8\��>0�0��
�:̦x��`|q-! $·!��̨DO���_�R	�{	9��eſq6��b��܀��w�q����Ԗ��{��r(���a� C���M�Bk��y��Q��T�Z[�l�0�*�l;M��ٕii~^(�HY��<����n�0 n��U���@M�6!��$�_{�#2�8Z󃺑2K����6�R-�S #�h��s׹��cNqJa�q��]�q��@�2�� 3�.�\!ݽW
����T��^l�����8::�2�]\����u*��L&>�;u�{��zX`�����P������Ͷ��x�;ف|�V$�@}�ڲMq,3ǥ�ӓ���<�t�f�TދU��{�Lu�6Z��Fl�щ�&y[��V�_]=?�+�
��v����p�i��{�+�M-�h�.j�{���}�9���bO���z`D*��
�6>p���҄���3����+k@M;Z̔+��E�4��J,6NP|J������H�_dѤM:���Í!�����w�QO�z�>[��OK���i-	鳜��m�!�!���Z0�L>�O���V�	neD����[��.��zM:��H��9���9��Ri1�a��"�Q�
�s��<.���"���CX'�觟��	e���#gjٞ�+)���S�b+�!������<�ċ�b��^���񇾢M�E& �]����5�4i-P���

�W;-�4�R����㴂�S��l=�+dvÚ���\s6��!����L% 4��[z&�����tL����3�9�x�n��Ά?*�ڣ{Ժ��m�d:���Sл<+|q�v�N���r�� �w99������5`@0��	���uf��[��޾'o�g-����J���tk�Gp�� -���w��㞊za�_ T B�YQU���1�������#b!�y�PT/�F�u�X�q)�O�:ء�٫���3��}���`�;Ƞ�=&�pyt�\�0T��:Sx�d5-�BTƫ����t$��C�W;H|�wX���qWXZ�9YwC#�%-��]�6�]j%�3_�a�tN�[�k����j��Uo������,��!`=I%і������j�%���72~P���!��s������䚏��6���gW?y�u��7�δ��·{��Sg�̺�׸�%���P��!6����:�$���I��e��#@��p�N-�Ly�$Bd���5e����bY�#�>m<G'CR�m#�g��c���������㽺}�G'�w�dkm���Kܤ�U$AK�n8���"w�[+�;y�3=k��(�W-0���� �#���oe{�$�z<38?��Lm���-	��NS����U��%?=;����D�Ϲ\,3�
�-@�Cf����
VŰ�`+�3-�g����Y�=Ʊt��2I&����1�)���v���[��
U�f�g����R��UK�vӝ�@B�߉���n�u���ȷF�O����$�e2u��i�E���|lu�̥��l��.B�q�
d��	�Hň�x��f�Q�6L/@��T�?�]�K d'�����M����7�Ĭ����g��Y�/��7҇�����N����Ú�S&��*6�!c�=�Sx���k��n3g>_AZK1��l�eee��R�Dg~��U`�Xw��P(Ɂ�˪ȍ����������ְZ�����
5�ڵƜ�Yjj�$	k���7��{\'����6�Lu�T����E�4�K&��r-{��B;�u9�{b���D�b�C�)!���sYw��Rpp�)Xጕh4u~�P��i��L����';Xv������.'vv��3j)��&�\�dL�����J�o�f�t���ʌe�p�f\+C�+R.^�(�B%�U9���KĨKgf�d0?�;�d%iD5g����x��vs>����|n�����L��ӕk���̀����!C��G>�
g�#O�o���y����H��ȺEp�{PA.�Q�`3�-��������[v5H�������9Q�Z.>��z~����J_�%A�!?�>ڨ��y|w������$6"�1C�r$c�|+��z0b-g�Mo_��ᴗ�o
��v��[�C���Y�[����u�'�HxWٿ*S{�e�){������L�Z+X� ��}��UF�s���J��[(�Q8"mӪ�x�x���D�K��*��������&d+o׮ɯ0�8�R�J�따��c!�4�8}?Ai�m�R�@���|y4'%��ج�'-�����7��ܙ��T���l���r�/�Sr��6K�h���-P�L����׏�x+�e�׺h�n����ߟ��_�ش��h���Ӫ�d66S��|�h���UWu;v�`�JEN6�zen?�>2�gP;��GI���j���X*1�\�w)�^���zJ�<m�;*�>�΃��!��j���St�L{x�LZ��i!�Al����x��	�r"��I9�D��^�V��O�r�)��5��e�c'���W�p,�WUcF�=� c@�	m9�`*�'��4����=���y��;�c8�[�;	p@ۇf�=���@�'���jԼ\�8�l����椯�F4�Xi��H[��2D���ɶ!m��W���2P�B�Ѷ�17v�����6orԵo®L,O�l|lTS��W���R^�~튁��bB�~�3U[$Q^���+Dw�!���P�)�nr�}�bJ��[y"wʵ_˫ ��&��uJ�i��h6񻑤�I2#=]���f����X�z[���h	i�s}�.������9��]΍���_���4^f�)���]��ݲ�azx�%����#��Tb�;x�ǜ�.�՞��<lc=�?9�9�$�Ͻ 5Gn;���ɭd�>aN+�Xf̼����x�"M�Vq3i�GRN�h�rg0��2Xs3N�-��A[H�M�e�Z�S��/Euh���H r��Q�ﱌ�ҺG���]���SXe>řU�;����9J���L ���Bg�+��c�9KwGtӍ�>��?�e2�2�"�@��L��]2F���3�|aO�r��$���T�N�C|�/Q�K�����E+�0�C[9�W�*1K/����匿A�B8�~v=���K��B=�r�����*l�"�K�3Y1�^A,��?�y�9��p������.ƅ�ac�-�|DmN}�8]�X:������q{�)x�v����v�ID��jh����!uO "ge�_�X!+�V)��a���㏺
��%��&��/��m���i�j�|�<�cFl^��cr4�vJ`��8�Kz�`�B1��׮54�[�� `��E���?�'������=��F)ͤhf8A*\u�jq�WR�˜;pȂI���Ս�BA�x<�N1�P!I�km��*M�6��D�8)e��U����K̂������~�vV�����:�4�\-���_��J�v�Y.�Spk���Yh��:~ퟠ��9���%x]�\o~W�	̊gW^��b���x���`T9���R~�q�W��)���Xx/���u7Gu�RP1��ؑ� �`�aG�������=Е5�Ѥ�	�'�=���v����d��߮Z�x��\�G��f�L�����֫ޯR�&�ʫ�M�`a�� �@��/���^��f��iv풽N�c�0G�U\�h�&����S%�G�`�M@���j�-oa�-�I$'7���ml�� 4��ɋD�w�`�׎�O������n�C
��~�,�WE�[;j~�d�۟\�r�ؚ�O(5�!���)��|dɇyti�V� �$f�p��
� Ɖ�WF�2V�L�����9֖tw����u�=���JK_� %��F�'�WF'�i�ǂ�/�$G"�N��ڝC9hAe���=A�/znQj{鷯T��$P}���Q��]���v�Gȫ��������0~�����.?�F&�v��
������ÞE�aM⋌}��@�җc��sW�h$h2Vn���g��ɇe�p@:_@�IV�]ܚ֩�<�TX���Zg�l��xU�7�-�����:��H�m��u�U��^	o�����^�D�dT��<Lt��_�8����͆�mKb/da~�@WA��[S7�N����J�x���#h����=��i?�~�@��m�]᫝��ߕ�<�,�����o��t_�k����$@��f�в2�0G��~���^�xnH�k�`���K��vO��rk&P��2��s��[�	+)u���c�"2Y�����.c�Õ��٩u���2�*(gj-��������O���cf��T��wN9i1���ŵ�Q���eH�^u��P�\>�z��!�><���R<$��M�vu�0R��Nt+Tp�v!���)��+2$m^;4J{�c�j3�C���j��Ĥ%p�)�;*��*n&����pOԮ6��lA�������=����ncG�E�٢G\�9[!!Æ��G/���N��<~,W��E�fșjqp��D1�u�������g���*˺ć�-��Mf����?	r���B��g�K�ea���1�Ty#�e�����_��o.�|�8��bg�(̅� �<���m�wvv�?:�ז����6��� �z2�51S���*7`�&�̼�BK���r�]��a�z��� Gm$*X�_S�zJ���6sҨ�f)F}��7/��-x��h^�+�:'����lA2��wb��ݞ�]|�M�9eß}&�u��w�G].�D��j|�4u/��y��_i�ߝ�;`ۃ�ڜ�II��zR�O�:��K^�UnT�:�������m�~�9\����$�ԕ��$"���p��Y(<[S뤓6���H�������w���yyIXwv�0X{��<2E���������jǉL	F7O%���*�Z�G��/�H��}�(���8�q�le��!�7ݣђ'�z�6 v�O�Hv�-\�����&���(�u= #�8�ࠗ�Čz�X��t{�$Q��E�[���`P_�^w}�h녕����s���҄CjF`�r���]�Mm�l�/,��9��B�iu�'�)v�7�\�+�����zqO|Su��u��B�`��L��ںك��Ml.;Nk��a�uϤe�=�~>��t5�Î�p�.�sqҥ>���<��h�����[ɂk=�R�:A9��FUņ�>$iE<��)�,_���IA^;�#��):���c��e`q�&�@j�.��'�&ar��Bi��[y�����s��+H���F��B�/�w����$t�K8g��L�����rW����۫��G���f�M�O^j����K�]o�S�_�o��ʭ����K�!�g<�E¶��Ⱦ�%�cr'��/ʯ*kE��G7���I�(#��2���l�|�Z�_VJ]�wt�V�W��T���;�LFH�<�U�(��i�z}۰�;��tir���fŽVQ}ݵ=��`QY,�g�M�W�̑Ά%�{��r@2@�r���&��6���)������؇����_Ժꍿ�b�n�b����9�H��W���W}�%��!�R7V��C���/@�������2y"�R��F�'��VŃ�t�3˟th�@����%���p�"#�b��o=��t��
K��fW��4ț��i��6Y6^#b�=p	;*:?�]�;C��]}�`mB���t�%ⳎS6l�F��%�Z*�5|�8��N�]��z�Y�o�\o������x�� ��b�U\�Z�w���3��K?���t����1d��E|�d4b�j�b�.���M2�1���8�<ha���^TU�/�
`�����#^�>ͣ8TX�*ג����K� �ێ,��/��$!Y�"I�!ʽB�Ъ���l%b�l%�Q����F)0%,����������- 13�7���|X1���^Ϯ����z���^I�=I�n�\��nU�2�~i����@@�VC�O~��&����@��0^d���w1�e�L=N-]��*?�0�ڪ7��艧c�"sT��'�a�wY�1a��^w����+��?(�G[��l%,�P��qmV���m�-��DWWך|���5�~/�՚���%9�Z���8҂��ۻĮ:K>�'Q�� ['(a�����������u��)�No���ɜ�
L�v]��ߔ���Z�K\?��@����q��U��۸�G�ѡ��.��;��rZc|��em��ж�1Q�R�O���u�؂�y�*W��Z��3�
aP�ڻbD�5����<:�_�G~;xϠ�e�ct�ϩ9�N��))��LA�mT�#��@�gW����xI�y�� ƂH9�U���}#�v6���שp��$���((�17ih8��B�E-����K_��,mVC	��
������k���.EA>�F�Kq1 wJ����\8�K3Bg��������p��|�'��j������ݣC�LGˤ��U����C�܀Yvd�����p�GO�L��y��,D%�UĊ3���쁼b����J�rL�--S��u<�t�=��m�{�v)^@�7��X�}0�z������hF"�Jkz϶��b*�N�]�X�������v���ݯ䇵j:]�b�0�L��h� �8���Id�����t��㒤6]��#���v,6������i�k�\�,}"h8��6a��d�k{�1��?t��������m���o������J��u�^YK����;���I��@2���I���>~��ΐ�*��^@�ˇ��
B Pd����Qypy*��Ip�j��6���7��t�r���Wx5�쑐}E���}@v���(XO���_�T�J[}_��Oz2h"HR@��.��>*ً� 7�Z��Z,	YK�$�2W`n���ɈJ�t�56���&I�B��]4�z����ᾭ�q�'vc��j����<7�T	+�=��^F(��s��i�p�pu��M ��w!�QC�%�{�(�ӏ5��Ǧ���%�-jĺ����~��>��J�;���=K�@^cč����I��g_�^���za	e�jwn��� �A�
�k�G�F]E�A�m��j�b��[e4��b��C�Οl���#���p(a�}g�$ ��6/���1�(mX�5��}����u�g��l�0�t��y��3Y�(o��|,`��������jqT�n�N��;�v�s�'�N#-���Q�m\͞�Im�]�ID��/�!P�{;��i�:�R3 ��������$Z-0�֯�X��Z���\�@��$z���u ;E�լ �m]M���F}bZ?LV�C=Ji�/�m�q���r�u���̈́���	*���0���
���4�?��j9�î�y�KU�2�uȗ��V,!�A��hxx[ʭ_ήqH�5�a
&q�ɇ���^������M'ܳ�}�T'�D�ԎI{&@������l/��G���a�WR�cPC���²N:�\�f�5��)e�n�\v[�ս�~�n_b}՛���W�Խ-��z-�}������`���3�"�J.m+4y惡����/`έ�@�D�
��X�B
��uԯ������)$ԅ��X�^w����#�<�I�Sꔾ��h� �B���)�.Qy"�F�Q���L�{t�ژ�G�]�I��`3stT�d�^�V�!�
�7��V��3��T�<<9
/��<LC�,��kr���'�Y��ܿ���ѕ��4B� ���,5΃@i��ūp-��bSh9�n���
�l�ԪNA�����2#9��e�M*����kX�n �2��`���nT䚽�c׸?��@&�QW�nǳ�Y��%]ʵV�=�4��ٕ\�k{�`M�o"o:x8�0y�eg�پ�2��Y��`�5/kMŒ&���B��p�?�sN!J"ꎐ��=Q���9O��]��s):�IB����\P܃67cU�E~gk��Ӛ+V�ϿdCK�+iTYl4���Aԅ�І�]:��}����+���㈆y		4��R���^�T����ǖ�d�Q-F����������3$�\��o�j-���.��\W�D%9�u�4x�n �ݰ��Rxtչ����E�� M�#L����R@d�B�r�k��5���J�2�OY�`M;#����#?!�o�x]�_��:2�@יv���ܓ�__E����v��[��E�O��2���z�܄��0\V��Mk�άap�9h�-_���c��m��F&�yl1K�XMIL���kuV� �rJ3���G�R8�YZ�m�< E�F��K}7�X|��af#�W�i��Z�Ɋ�/6� wsf���w�kP�W�Q�f��0�9��=���h�eH��Q~�%�����ǵ>�7�Ӽg-�<��BB�.G|:y{�޶���p\��P"�d��~Z�,�z��ե#E/V����s�v�M�5D��"o�N��a�;v��}����~3S�n���{�X
[�Æ}_eu����Vy���.����TH>�=��r.��t�ut��W~(bX	p���|S�u�FH/iL�/��a��-��?�E�eY��&���d֎��Y@��a�K�0��{�uF��Y�����R����2���H0]/�c���*6���	̴�������������n M�2�O3߄��Bl�2�n��k\��vp�-z�~_�>)*����)��I��[��'�߷軧x�?�y���g/���wMVA�v]2Èg*u��.����6F���3�W����+$j�mWrR�[	gpq	�F߹�O]�[м�"K~8�|�.�:c?M�]J�9-<��7�R�kZ���l����DK����s��1��佴�*��v�ϲ�8�1�ͅ�g� -���<����7�2f\�هQk�F�M֡F�U��F�S*
P�d��I�V��|�J��i返���@�ؐ+f��^#1&4%�;�ŝۛ��1@a1k�vV�G�b��݉�wGR�>F�F\h,���R,�>F 1����ja�����o����͜��0��D�&��0������6Y!j[�dP�#�sV[)��i���`�x�b�����P�Xr\�/��谖��G��3|5�_��{QONn�, �K�d�+�˶�M�)��L�7��b�S1?~��@�o	����m�ҷf] ���J�o����H|�19\x�ڜ��5_���*��IQSS[�~\���W��)��Q�������o���I��O�*��R\T����E٨\Z;	;��3q	��*��q��Xѩ��xB�x�>�sq�B��o��}��{N��+I<��#�+s ~wz;�>�����T1�~��bf������کj���ZC?���^���j�.������	��S0O���G��*��\]u]�U�MJ 36=���IK���Y��a�Sj�Ϙ@�L��	��Q��7�'���Θ�"���l�� D��(n����3RY�����l=S�%7�k���X���2L�@��X%�;"��"$l?��0d��
$V�۲��t���\�V���yTlo�%D����� ��D����m��R��!lg���lz�����}��U���>�	�9W��.����<��� P3�g������Z�a�*J�F���n�K���gq�m�aX�����T�����c���4W����j+_��I��#���x�6w彣�����W�c�m��ū��<ϰ㬨�t�\;��W����@�r*�
2������#Zؔ��[���Ԧ^B^��[�V����Wq����N}�I˛��d:)Ǭ������RD/-��6T;��p�ro�nsm$YE(@AD��ob���ͺ�`[��ؗ�& c/!0(4����f�&	,E 	)�{y�X���	3�OU}����`�V$vGtjk[�[�.�Q�s��B�MhL*��W�pr*���3�k���𯆀���;�\�y�����_f�Y�3l&@���_+d齎-H��3�2q�iA����q�]�9J�V��#�@�r�\��DjuݑV���WZ�[�b�$g��J�I���aO2��<��F�||�I#�T�Z;�x�����`�zP3Y/����1b��D��;��&�dC��9�W�<�V�󍾆ZH�w��ƨ��<I�~��,)��Ҍ�8%:[+5<�g�6�u��5_8��)::��Q� ����?D������C��m���]��s�^�^k2�@�-�i���$��x�g��CB�U@(��29�W��;�;o4q�V�m��$�y��i{�ٻ�����{s�YCm�'�5&�7�)�;6���L$6�ܑ�����d��UH��'�A�Z,���n��iF�ݖ'��|)��`�x�$*�u�?__��x�'�n��Wq`��$�(��Cxk�<�\�6�������w���O�Ņ�e�ЙyL&�>�3_��� t�.w�g(���z�-z ��>c)q�}��YL��ǏN�P����U���Ɏ�[5�5H�d����j���0F�Hw��xRb\��6`R����h�����m,���d�a���7�t�؎qCn���e��=�b˵ä 2�BU��[7�"p��g�'S��zo0}W���eI'�LS,�Zܻ����8������A��p�#�|.f�2���ñ�r��5�u9�3}�M���3�|���X��̵��n�Zv��g(ǔ�]͚K;��V{2.(��F���镵��%�0�nR���LǕ�a�H����=*�V�?9y�������?�a{r#*�:�!��'J���H�А����׌T@�y��
����ٛ�<�Y\'����-�F]�r�?i��~�?A0�/��멡�!���KW��t��d�K-�o�Ʊ���Ά��lSQ�k��n�E�I�J�BB���:|�^��=� �D��J%H�S�(�Y�*p�Hfq��`��z��{��n�Yl�MT</<|��I����5dt��ﰇu/^*B��Dnǚ��[T���p�,n�koP�
��[�Q8D�����p-�qV��vyO�}����v��E���o�
��S@a�;���[�3Ln]�p1�Y�Yt|��[�7
�����ɤXI`�w�Ĝ�#_���tb1 ����|�NU�Rp���9�qo�����O����E�D�+��!�?�ޒ|<Ϡ*�d�dm�#��!���-y�\�?ފ�F4�S���&e.������D|G�Ą�M ���S����Ы�����{d	��a
O�����	��F�Yy���@aA���k�9�m\F�KW���z�%#)����9�R�XF�^l��t�E�����Tm��d�|���@7qЭ���U2�A��u����2O.�mNտϔ9�v��U�q"֊(��Ξ��/�[� �"��ٴc�"�Ȼ��t��� 1�l�bs���/\9��kN��BH�%���.�J2�\��i�q!�4/*y���W`��]j����_��>{��pd����g�+���tC_�Em��X�W��&uAA�W���ɓwR,��R����L�R!�)cQV�| ���$�] ��T4xo粰j?�����݅3ʕ�Yǩz?����.�ru��$�=����]r�ѸGmPl�b�*�f
fN/�v*�#��m��Sx�\�p���3uL��$jkA%���ע�� ���;+�wA�V� �<�=hU!oX�EF�;�2|8���	J&�������yL�a4����wE8�N9�B�2G�@8�<�Ը���u���/�z7 � �4�Y�&��{i�b�B�|�XN�cÑ�	��^�	�g��F�tJ^�
�ѹٱ�Z����[�Q6��>2.�od�����,W�r�{�C�����t��:5OO.����_R�ޝ��x�޳<��D�S~�9��AJ㺷w#^	|�P�ՠ���<)�E�H���x�S^�2�v�b��lW/�V��rK������E�u's�d�_��eٵ\����4-����x��Q�	�һ�C�C�{�"����S�Ao�����<O�3�]o�-��w���7�r;.$2�O`W�A�-H���������-?���"�#��	W���8楙�̉{����OyQ�Rn\�����4o���5�j�b3zu����u�D�9���PEa�b�2�3C��Jjb�^7�|w�/�(S��de�$�{�^c=Pg�Q��c�ys��I� G`��\y�9����3�\g�%�^T��ܫ ��u!}� 0��37�=0���p2m�~+��n-1��KT��=�a'�FP\-�v�pZi1��pt����j����7�b���������"����x���j_��!h(]��3O�D�F�O��f������{7;(8�w���ȍ�����'� ����Fr�&�H�����#��k�=2��rb3�����|���G������]:f��0Z�)�-ve�2��*Y�ŐCѾt���b��f.�/rk��}lN�]�Ȱ�l�˻�2I�wi��z&c :x�H2eW^x�+���p���.���.�_K��������ۋ0��|��}��
��u���>�)1����/�QO��@w*�Aު����Fd~7BV�4�گ����*=�6�Ƹ"^x��ǻ2w{���{���r/���m�W�9��ӎ�[�G�Ӭ�Po5 �����Q^;,�<�;�7#j�$�#�Ck���L��r��[F� ��Q��.��z������j# ����� ��DRnw�k'N�F �'�UA��.>���.Øn��eo^�ɓi`Fm��?�o�Hw��&� ��~��y���:8�V|N
�d�ȯӲao����}�&e�Q���]!�5@�[@Ω��"��b%���}K��Y>��˿�`�[�2�9�2Yh�I�W�"�Dޓ_%�5(y�<�޿�"���k���H���j�0��e�V�[q�&�ʣ���k��T�JL����q���X���gUd6�uGj@�W�{�0穡-�������t�Ɲ���ُb�p�֤tDѼ�},�J��nT�6��Y˂�<=D����ً�4�"`��a>�ǔ�T䢀v��ϼ���6���FQC�o ��_�L�<����F,���O����) �y��y[ R���C�=��[���W8=�VE����W�5�vac *e!�� ����n&��c�0T�{���ݠ"  9z��c�t���=����}�|�����\��+@��}�	�،�� ������9�V��������/,��i
/-9�̚�������sMhL��QR?i�2"���<�e��>���;�/�VH��,E�U�c^�ΫA�.��W��O��ԩg�F[�{[�xVh�`Y�>
�]�����%��GXk�]�2�//�~{�S
	�{]$x�e�X�|��y���^��!����oa��˹�	�^�?e��5ݰ5x��|���ʹ#WS�\jU�p�i�"�=�"⺎v�`Q�N|0/u�ad�}j���/�l�~�HBm�bu��n��&� ����lo�� r�+�	��w�_\��IS�e�z>�A�֖ B_$P[ڠ ��@�6J��|uc����?�5X?���X!�$��˚I�l��AM���k�)3y_�#l��{[v׸;Ao3f��;;��ٶ��|�^IPs1�\͓�H��k\�Z�cU���[��!��4��lqB�_�� ��P������;��Ϸ�j���ګ6_���[�_�(g���A[�vKVl��Nz��g(�릋Lm���%����bD�I����g=YsL#�\�,�l=ȱ����J������6�9��ܣ,������sq�r &`� ��4+��\ӳ�F�q2��U��m\���B�۟?��r~�dKW�jBb�Qj��򃶻��tr�I�WT@@JL�|>ب?\#�{�X��6? n�F�$��f;��� ��������d�����=�{�#OWv4��D	"���γ��nG� à�6��o��3���=F�$3��\��[/��	_�U:��Ơ`���G��9K۔'a���#=�=xA���j�eJ��~� :���&��+�=�����'�W"��Y����Qx��Vٗ�<�o@�rO���@��$`����c��L������v,f�o�>���":�}y@��m�����癁m!4nD�je�4�O<�����PN����e��B5�z?!�d,TSdwHNV���pF�Q�{���t���u9��a;΃:���X��RR]S�\��A �?{u��2��{�������\e���wx)���:��5��HH�xC}U<W⻗#˶; ��[|,�����9ZȔH�r���������X;0����R���7��;��9�e$d��>��ޡ����o�c9���& XP?G��9�H��bqt���3=/�2�[N�3.G��Cl�w4O��8���"G�5^�]<[�#���9����֤`�a�/�����t���彔��°u���ް��(,����鬵���1�7�3�j��,��~δ�:��R˕r�(��J���\�ǈ��v3��/K��a����FN�w�χ��:�{-L������!f�srC�֪�ߕZ	Tگ��7�O���~�Ё
n�Л����� ����?KI���1S0l.Lt=@��Y�� �QF�?]��E㺦��n����t�v�nxn'�-�y������"�|���w^;�GGof�g�f��3�Ys�ٹvv���l���dL�d@��5�aIپb�_m�wg�`:i[�}� h���Yv�5����zx���Y ��l�Pf䦦���ݥ�Rx����{���s��sn�}��rc��yO���}�hs�S�E���%W�ўOv	�H��,�4����{{9�X�{)/G�g9����amQ�иe�{�Æ����Ꮃ�v�ߏU�D9�J�^�Hdl��B�8��ˀ@$k������b��5]a������O(���q�T	�i�vLIiI��T	s�T_;�
��~�|e;K~�!$��d���s�������s��.��y.���zAe�M7�=T՛�O��~�����
w�f���ɨ{^3R2�+��
+�	��I	"JZP����9��rg���2����mN��3JՋ/�n�g���5��GT�0}�п\&�"��8׈	�;�E8�f�Oq;��^���
A\��]pq���^c��σ	��/�̖���Om��2u>�oT�_���v� ���)]�p���nn>M['�� !��!+�l^��ъy#�~Y~��gw(j��8
��I����!f?$���\aÏ�*�ru
�vvV*щ��Q���0PPK��CʭO��P���K�w�Ú�� ��-�Z��G>j���	�)+�������Cju:�	��aA"�l7�^Z*"���V��w',c���b���_�:�������U��n���˻��N�k'h|/�G�\�F�"�2��!9��O����*"\;�'��eh��ؚ�GE�X���W��r��;�VW�UlUZbt�dEbQ9n����{��R>�_�
�#ٱ��'�	��؆_��gpG�ǯG��'G��:j��cj���4R���I��'c�J �K�>��Mٝ���j��y�I�e�7o�b%�K+r��.�n�4���9̘~����иE<�[��ą?��Bs>;�A���(�#��ݧ��!O�����-@g�d�Bn����4��H�;-]�{�������=��� Λ��E�F�8�aOާŰ����v��#�ꗃ��]Zc�:�k4�P�a�Ms����VC�����S*'+g������x�b_�l��������pFP�]/	:d�-x�F>g��!E������1A(/��Ѡ���#�L��A6�թ���ڼρ��wD�S�� Wԍ)Vf�Pܢ*��[��v�R3���������6u�#�V:�o?��P@�j��!��j�՟�5�7	�ڴL���<�!J.r&���|\�y�	�'g�vhu�R,��K��g�kN������J��J�d�Y�.��/��;z�w`t�b���R��`�P�E
�]l��9�Ӂq탮�,����*!�'�� �O������!�C�Y��(�m���q�����	��"f�_��L
d�Ch�����g{�oVV��"�0��z!����i��;5������&r�զy�OTy�d��b'zuc8�:�<Rc�F�A�A�j�4~����9*��[��VH�N#L��j(�MӽM��K�rm�Ӏ�Ms=��|��DF�)&�"��ϕi�6
6�E`
f��[��R/�D�մ2DI��ߪ�db�������;6�ލw���.vdaS:d�P+|	��YɃF��R�cO�4��9&)��4)��v����7�	?7�JR���>PNy�O1�[�^nog�ɷ��t%� $}n;��{��(\B�҈n��8`Y=1�۟㝡Wa�MO5_����]��2Z�w�������`��\�Ʊ�鐑�a�i�J��0���$��N~t��g>"��~�����T1a�h��}\�4�S�>�������3r�m��*�OA&_�iq>x!g���%Q/�u�ؔ�Cx��a%�����ira�2.YAS^�U�l�?���V[�'�~|����F�C�����,մ�U�W�7s��>���{Mi��5Z�:�=}��m�0���莙��ߊ�Y�e�6D���әq���ݩ]A1�e��i�e����&=��lmn�5�KU�3.��8O�2�' cU'����oU?l�G9��!��Y�D/Rs�ot�N�y��۟���^�6��L&ߨ�֋���YG���ˀ+�{��9ޅ����O���,�|D!����˥�^�~�Qn�)*��\�CY�8O�/\ԃ)K2 �����1_�R����g���7�����\��M�vZ�JJ��j߷��
������x�@�W�٢G�����*��{h5#%�fͫ���&!���;�0��{��T���F�Jځ��qp�ßc�&M[�k�Ӎ�0Cvy*�I&&�u�_�m�'�ήW����������buJ�}�D�Vݶ+9�A�En@��y�:]T��DXE̻�RFj:!Xt�4����z��|aGC�������
w*��t�N����$���ɜ��f̶��� �O�j�-����rSE��oc|`�9[� �?���v�*�Ѳ݁�6���Z"x%����߳ T����"_���|��9L��a_i�e�Z�&e�aXUq�8[�p�����M�z�-Q�䔪g�go���j`�Q4����������oh��t���w�Fv0�����3���tHu�)�$]��"�\�m{�Ź^_='F��R}(�A��et�J^��)��oW꿘4)�@��q6G�[��ʮ�&�	���o*;m�V،%�^�iB�o��y)�1@l]v |'8��gs�����{�;5e���ea�!$��Tb�t�b?aF��W3�V�]D$���R2f��x�Ú�ml���������>�T"2.�����Hc�$D����}��
�z���l�k�@%�����a�,3���D/�x�|=D���&nڋi�:6Ǧt�Ҋ?[-j����ۖb�'�2���	�]塳;��}�;��:'�k�L��!�[�
��$��>�?�_�=�ٌ�;����ML,>�����1�|�W^�KN�	��+��e�
�E/�̀$�3$�*�y��׋��9ާI�g߸:���������r=2�a�oe'm�g$�t]C/Ul�h��48/��T�>����d���$�(�y�yvQk~ş=��2A���v c��?��?�j�O �:Z�ތ�:	�s4�Fl��q�����G�>*��Ns���7�v\څƵ++h��J;�'��wΆil�_I�O{e�MĊ�Kr�6�����#���^L��g�&���,e_��b�%o&F{9�z��O��+�a̰�q�}�r	�������~��/)\˒���ɞ�Ϛya�n����񭰍m��}��)\����%�&����a��g�w|��\�)�L���;w���z��|Ϻ����n@�ȺՏ�fvzҳX����V�CI��=Z̠��)Si�$�W	C�ɿ�?`�ۘ��.s({ob ���c����E�����m���w0��@�;�@k�x$ָ"�Xa�i�R,ee<0>��%�l|�yw
B�s�Z�=|���W�Pۉ��Y��ɿ�3L����3ū��N������vP���'����6�kT���uYeM��O�K_�ޕVn@>�z�uMc�)V�38_�N��t�Y�.F�p1��
#kbފ���{�-����x���>vw�H� $���QU�T4��>�����x^-���?&／nЭ�� ��&6j����S���\�������d�<�F~������4��e�����9��ƐC�奴�]�AJ�|��nۑ*��}�_�S�K�X0oYV%�35���&lJ8\�J�݁�w}Ao��
L�� ]����u�fx�o�P☺�����j��44�@ڕ4٧ݩ"�3૦8F˧>��E�|��� \��V����+�*5\mٸ�o�fg�`R�}}���B*0���+�O��n�pN��e��rb@��u����KgT�} �o􎊀Y�E�l���es���I��)]6�P�PY6�SxS���L��Л�����o~�x1��O<@�{��ߥ���"}1LJhB����"z�#�c� 
�{�|�e��uh��e\�FA��O,�n�=�?��ܵ阬!_�mtn$��.�QDuX��B�j+�o�{O�Ǚh�V���(�V��b�b��K�p&�J�5g�
��(.Gϝ�,�]e�� \�v"N��[g\כq��G���2�
��+�U�o�b�����ة�a��S���Gϓ�ZA�K}B�A�lw��Lp{k" ��@ᭆ�I��f��C�
H���ˠ��'ֆ����IܶwIF�@V�����6<c��7:�������(�������:����Gg�Oܓ/��ɶ��cb�h|��x�>r����Փb��+e�P����#�d�i��=?�s�(�v��]������o������h����W�z�t��P�`Q_�����/�޼�#�wl��*���5N��f*�RA���c��\Yo�3U�q��U�(hY����յ]z���1�
���&�+��ԃ�#"}�i���Wl۾u�s���[t�{�5�8W���)7����J����΄kjǩ�%R����Zi���j�%*��f��y��?)�n��:)=�]�>e䤫��.�N���1V�=�x�t�i�2�)�S4�04x�hԾ��`?�XoNG-�Tݍ)�����V���ՊnC�#�V��ķܼEk
�0��q����xF�U&�H���N��u [f��zK_G�Z�ڮy�zEd0#U�Z֠�K�oe	�f��lr�����9��@�;�k���1qL{��FL���������g���#.�Y��2������g# p )�&U�ht�t�ns� ���wِ�+�٧�o�j��!)�l���G�F�>��o[�+RQQɔ�hj���hw�Ym@t������޺g�}���qZ��
N��7b��O�Z�������,�FXW:J6�AB'�{���j�@p��}�U7_�.�U���Y��^�p~��5����`�#�nm^�J�\�\�^K�B�zs(�����w��K���yJ��>=��ʅ����
:��m���N��:o��Iz�"B�b\.{,٪7ҽ��w�\�	���5����tQ�Ȫ̬�+M��0\�'�TE��[��M�-��~R����9�2V��$�\w�nq���q�v>�����y˪zz��K_�]�g��'S�̶�M�NJ�3��4� �ͪ�OR�Tͬ�����L�Y�W�a�e�M��֔W������Z$���
�
����O�/b�]��\����77�JL|�\q(y�Q���K���t�V�6�Ě,L�{���T�M��M;���.�	qsJ�"��O�9���^�|D���oט��<c�|��t܍�I��8>�h�U�U����uLl7��ѓ��3i��E�C@�qC��7y%TнmO�f|�}��K���lƮ�	��DDQS�&� 
����v�R�5�~���)�bu�������T���'?���9��~�#��į��/}f�@:�-did�[8�.!����]G����߱(����Ր�(�>�I������EO�h�lI+�fz�T��K�V�?}j�ZJ�� ��{E�b��ӈ]L�����ֱ݈3w��N�u���h���V�,	�H�b˼�-d�gHe%�l%�)ò׈���������E��L�cJW��U��K
s�tlygggtor�?��XNDAl����F'���_���|�A-c�c�;T�k�p��J057'0��מ^�����qF4�n����Z�gx��,�ƲQ�bSvH�r	/o2~-��t��%�>dӹ��i�����^�b1��*�v���VӔx�\���d Ӂ�������$�'lm}c��saIT9DL�	h�*�77�#q�����r��-GS�����N�z�n����3�����1�v�E�G�sU������(����w�5G���{o�����^{X�ܷ`�MOΩ���$ w�Nx��wI�egI�T白�+	�P���u��<ʋ�x�1���VV,b�r��wtX��0<��G������^_S�af)��Y�<�����E_`^��J��6@��v�k4��,�F^���n���� �?��mCEA�2�N45Vc]�%���N�Q�*&3K��?3��������>��1�(}���n*�6*�c!����t�\e��k���D��^2����=Y�t���"�oRVO�CB�p�����l�����*�V9���^Ot�̪Kq��7C[�OF�D)˳��*:�E���cRߘ�
+ɝ���>�hxN�Io�?�L�p��'�硂X��N ����T~o�s��&��ț���)M^kȰd�i��W������ޯ��W&�X�yi�sy)L�.a�Y�պ�;m|'p5��"*G��4�޴-"�K�q"�����a����W�X�SU)F���������(Ժ�u�@��6�/�$yZ��_J=|1M�qp��Ūz�����^-G]���8A���V(�� /Y���*��N�����ʲ�Z�_Q�1��"w������E-��ŲgW�A4a�ّ�se"���[cK!.��m��Uv�~�eֶӮ׈-ߣn<_�Ԋ�}�w�&�Z��ƘVޞǜ�l�n��l��.�H$���|Ԍ��6q_h����g��Ɲc:
+���\�aE�Sxfu�����w��i��Y����3dy��@ ��ly�n^��ai"#�6��}����N�d��!]2i:�ĭ*�ng��醇�:N�,igrfr,���u?oʹ�������=�85m��P����o,hZ^Ӵ@ӫ<��4����=�`���_�Ϧ������O��1Ѯ�꾘ir�����\��O����ߖu֨����i����_}�3تbFg�ɏ���/2ɨ�� �C7����xiz���o�3���[����Y�6����Uq��)�U /0;4��m�O/�..�L��b�6
>R
f�}1M����q�=FHsj��'Dt�͛A��`�3��������z���9���H�C���)�� (�6�B���m��ھ4R9~�M�ylO�h�6���4lh��ms)��Tm�z�I�$�}�G�0������A�Ұ�br�I�4�/�wvj�5Zxly��?�=n�E�Qj�8��~�g&%�8���SOI����,j�/��Դ�M�k��h���t6r	{��?T/�կ�/k(i�V|4�t���qx���4���a��X�/[�ko�
����C݊���!�����x8����A?�{�y��y�� ���^�G��d6T|�f��c�����pt��;���j�07'��C���٢i�Į�Wv��QC�٪	�c�W�͉i���I!�}e2�{+�EL���B<Z�j�e��]L�^�,��zw�:ܽk�cZ�%�핮-'������[�h�n�SuCnB�o�j>֑s����،�Rv[U�����>�V�b��-/,y�?Ø�z��f羥a^�rÙM;�/5��W�Ж�	<�>f-9a�~v.��&,�Es� W��1�������x< ��&�)F�P����i�*N"���p��<�\BB�n��p �ԮaM��w�cf��&���4���=>��?O�V�T)��A� ����;@�DN1�kF��Ʉ��$���� 6 /vH��G�V�;�����s�;g]Q����L��w]� kW	�Q�D4& ���`]�Ԗ��=��t;��έ�y_�~�ݺ��c���c_���hY0�K�"���H�Elʝu�c��z���#}b:+H�/C�?��a�r}W	��>U��݄�jS����|�"�~��|�?t�{��E�����q��u��t��|fUZ�Tσ��u~'����^ x��\�@2K�������+ ������n�8>�|�dP��:��f9ejX�

Sܭ�U(�j���͛�Q��G��M����&�#��.��]5���['��$,�_�a�I�F$�����۫�c�XWM���Y�j�1��"��K�.�^���@X�߽�C/27��kc9�l:��e�s��(��P3���{�}��٣���g?Q�
'U��1�m��\�{6�ҕ7�=P��:�N�51ǪX:O���Ku���%Y�츍\ ,�:r��5H�iJ`\_z;\ޫ�H(+����s&I
y�(����q��{��r���SS<�K��TS���?c]�ö�zWPLW��B�x�J���8�$vs�}=q\�1ӛ��g։��m�5�.r?d(���}���x�/^�ԕ,�.{��_���b`�q�����a�J��8A�����mk�`���7Uɋ�a �Ș��a��l9�=w~ϙI_�#�I6���뭬j�"5���z�5Z��ZWY�@�d �Ķ���7ih�%�"2H�#`����C@�9�=�nm��v�4�F'��̙[|��>vB�xM�f��&
�t�<1>�rHl���Ŝ�������m��FgKp�~�"Zm��{�l�-v�e�}��/%���n�H�s�I�~HuR=��ӷi>@g�^As�^*��	*ϟ���	b8��/�fVw<�e��=�b��z �����ķE@ߟ�**n�e�ZNLVҿX�ݷ� r{ ة���H%��씌0�^���E�����У�%׿�Wڰ�:-���l�����Y����h
�4r_N����ϛ[����ʋ#�;Х���<�F�.�ܜ�OM�]E��[���}y��TP����Ĳ�9�K�_	="R5ap���R��&���y�qi��Y��n/��F��у�s��G0��Dye�e�[��TMqd[���V���+��D<-@\��(��Id�&N��.�B��j��]ʚ����-cs=��Mn�i[?�o�Mȷ۱2a�\y������rJ�^���3���m��AQ["򗂧��?��A�T�T���{�S�0�Ŋժ�w�啠X�Wv�Q�wZ�r�Ne-�b0���!W�����?;}lmfc15��o����Lѯ6�"���`<��VT]��L}M��T*���4�w�_~������.��Cֽ���1�R�nndU�G�0�1'�i.x�Y�*��~._�hW=��.�=�P�ˢ�;���E��8ܑx�A6�V А�	��{x��4����>g4�	�]\.-�\{��Dɭ�
�=�D�;N(��ڞ���B=��+5�����ީ�_��*b���iG��Wl���D�z-2�d�>`H�$�#!)�!4vQQ����������oܘu0�p��B'�4���4+U��w?X��6�����|g~�|�����g	����w��kI�(��q��i%�b���D��q��O5�U�%��0%��Xqu���-زq�61����O5-�fi����k��'�P��g'�ce�׃.�S;eI3�MO�f�g�����n�i����p�SRmj%O-G4�������Zhc{�>j0���D��e�rѦ�v��9��Dp��
Mo��yO�WF��#6�j(Six[�����M��׼��$� �*{�UPI�l�@_lw��[�5\BD�8�A��h�֐@;un�~�.�C ��@(!.	�	E�.v��e.64W���.QQ�-��\�0�O�Ą��|��Y�gFS�4���d_>��	�E���v�D���N�q�?k��ɱ��K�]O&6������D���<
�L�٣��.[�������c~À}U$���e�C��#�z�j�)�M� �6��~	|���'l}2^%v�zRҮ��Y��?9�#z�7^�P#r�J��ޯ_��:���s��?
�X�'�j�Z;`9����+���Tl�m��Nf�����ax��K���>��1�n�)���L�A-/���,��l��, Jf�z��{�"���jTe���fKZ�~��q�2�_i���R��}�4�'����"PPX}�O*4��x���T���H���DnF���~'n�B���A���� F�e����C�	Ա�6���
�~>���rF�٧P'Hמh�qs��W1*����[�������w�0�}N؟�C�|{ҥ�ŏ�[Y�[���gz%U�꥘��z�$�T�f�:�ɗF%8�cVɔ���`y��ٱG�[�{CkUش��'���ɟ{�1'��mJ1��9aͪ��B�Ͱ�"M��zI��4�Ų�v5�+}>�`X��d��M���8W^49b�Ӫ���p��Z����U��ۣ�5�Ϋ~��g{$����'s�S��
�r�ʵ����1��})�K�K���Ʈ �Q�ROX$��ʿgC6��ٶ��i�3�l��O��7���=X0jQ_Ѡ�����MUx6�����|���X&^H́7�
�L��D�Mr���V[�QX��
b7�5.df�kU����M�S?�X�'�G�t旲J���gR�3�>WO1�Q�szȘ��u��-�J?�ke�)��?ԗé�?3:��IIQYNwH�H����������������U#�5�K���]h>���#<i�Y�"�S�d�5�,����7:��AF��ӓ�^�����p�m���fYj���Kϣ�+�C5>��jW��պb%��/EOic�.�R�B[A5���3���
3b����ձgKB��r!G�����<u���.�]I���W���jE�k�._X�`�3�H���IL�B��b.��*�B��A�O1ș��~�vc��p�̏�-l�$�Ke�e_�jR�#Y��\l槬H�4�צ|�#��[#5��Q������4�&��(f-�\d;WੌY�Q�Q<n��Mml�+)���p��u�|h�[٫A�x�@��DٿX2''��ӓ�f2���_N-��`㕟��*��[,���=9h��C��J���F��:P0�M�����������`�@B�S��@}ųFܗ@�JX��o����%T�%
�8nI����.�J�9O���&��cփ[�;g��\�7�au�����&kb��U�����`���D�&�P|�NL��Р��C,���e]�*���.�5[������v
���}���lmR�͛vR�X�"V���u�;�IB��/%<���.�_O�(
w=�LyU���Ù�\<W[�1�	���&���#�&E���ĉ���N�s2��-�1Q�`�Y� ����pi�V�G
�z����r�mte;��вԍ@���V��SUwᏦn+��s�{q$w~�o
���u��A2��֧��Y�^Н��)�"W�6M���W3�X�u�i`����Ŕ�%�����\qlX��P���YhFV[:�s4��.� o�nv'��iy'�8��Np����ɧ�<�����<� ���w#$Ď���D�y��+�+�["�8<�>b*ğ��UΜϟ��(���2
��i���bwr
�m`���c�}�2��
2����@銕:m��C,�g3�{{u�����q,1t������I��"�h7��̺���_Q*��6��c*g�oȵ��i�(�V���۵�A�gx<K|����ܶq����N�������\�ӭ��W~P���2b�A�Щ���b��ѷ�&��(�Ri���5j'뻝�����JT�z#�, ����;
��p4Փ�r�|5�7� ")�C��K�H�PNt�l슦�z�
hB�����o
Ym ��V��]�^�x��_��l��&�x&E�l�j�$����{��k��G���z��������%�\&�T����;j���������?6����fRN�Q��S1G�1oq"�ĲX;	a��_(2�Vd�<ۍ�Ze�?A�}�\7�}��lH�iG����QD��X�yFG�K�ǀB ��BЗ�����S���h�WK�_t �C��!���G�E��ޖJ�O��o{�������z^�Kc�4"KfI����������H!��b�m��ub@�jh�&��Y�ڕ���-�����{�޸�]{$�H�@��`<�
��T��͌|ۘ�}�i������]�q�R��p������F��\C�����LB�ȚܔZ"�B�#�ƃ^�Iܨ*/��SE���r$g��f�M��F�mMD0y9��$�݁�OJw�� �#���*��.������
�՚5d�;w�I�7| ���`qj�$�܌q[�%��Bt�?��*,�"a<��^����5g������<�ug%r]
����Ҧ���z�l�nl���Z�Ը35���Xl�����[.i왙�f3�� ��˾9u���>(3���1�ٍT(Tء�T�s���oSB�~�ӊ����Ѥ]��΍�=,//���3+�F3��9o6-���w�{�����]/��K2�����܇L�7�A	�x��I�K%ץ�1\]�D�H�&-��*����O0+nl�"4����1f"2ۦ׳3˵������M����[ٯ[���_�+����]}�B�y��!x�c :����
6���-9��aY<GR!*2��q���e�E��Vc�Q^9�?B��w�4��mȥ���!�tu�<�U�[��Wײ�_]Ӆn#x���0:Kã�r��i���[��+��癔�0�=HUs�E�	QP�ӹ��E(���^d��D�iU����k�{�� {�?i�|ÊP���a��yZa��4)�#m2˱��ƉMk.���־�Z�<N�{LꞱ/��,/����X]�[�,��/�6`���'C�|al�_��=������D���@;��C��i�!´s���t@�����mJJ.�׼�bz%^�YNg�t�����9#H��G��(�)��(y�S�ӿ;o�yQ�[ Kba�*�8���5�����\����O�3,�kP�-F���1v����ܕ��4��K�=����$���iNK����+%v���n4���+۔䜄������f�{~��J�!I>��d�=�M��'�^�e�yx�Nu����<���1�_C�����}��956**�����~{g���v�m�¨��Ն`��ZO���ىD"������
~Mq�n�q޳�o�`
��S܂�'�->�y�%�L��_5�3�����>##C�)��R�Ѳ�>:&f4��Cِ�"�&�z���b�pggg>Hc0��ʋ/X?���6�����_i���������0��0�p%�w �v���C.����?<�������W����ꥩi���x.~��]���3���\�-����F�U��X0��^W����r]P���G.<S��ݙ(нqd�PO�K���"�"��+gv�����w1		0���D
�f��.IvEf�$��#��{�������J��ûFϟ�W^dLv�q5�QRZ*�
��Y����7��,0bk�0Le��FGg��)�0�lwr��v���.�wFrE�E�M� ��0�G��;���y[��1���+�c��+�44\��p�h�3[A��aj_�z�V���Bz��57��~�6�c�	�>55o߿�Hy��B�"���K�[\6�i/�������`'��U��E� �?�Q��ty�4W����{,R��'�ˢxg ����{���	�JJ��������V�����bӀ;�_C%����rT��#ݾY(e�؎A^ߍH�B�|
��[4���A�R^\5H����!�s�=�̔�����w3��W�.%��OY<���6LNA��u�,!�[p-���?ن�U�t�D�w|g���Or�[���ڲU�^�N+h8���hg�/��<a�ׯ�������E��[m�.�?	��A�� ��ۈ��y��?9麿!g�EWR�f�c�	X<)Ĭ-��t�h���V����rz����0�/Lth	Wwo��A1>��s�䉡�&&�������-)��0N%=�|o}�Ts��{[�H7�)����o"R꯲>���Z���Cn���y���z-�DEG�B��^}#���H�,A��Yv�;�ۤ�
ȕ�A��̕�HM��
��ͤ��O�A�
\�n7��H
����$u��K���$a0o��c���c��U/�8�c ����[��H"�ߘ.{��N�Ĝ��J�e��ћX|b�}g2��:�_�tZ����7�}r�2�C�~v7o��Y�����	��s���Ň�zol�,�Z�q}RȆ�5��W�/ffd:7t����l	���kx�Myw�N�&�w�����I�_A�\����a�V�S�߯)���%Z~kM�5��p6�6CF��ޕ���.��//+��ɑ�m���)�˫Y[#����k� ����c{w7�|HF#����BX>���A2���5'Ǉщ�}eu�
��y8� ���, �?k)(|������r����505�p��Z�b��}8$!�k��1yR ���z�� � ��^5g��V��/�eZ����' ����]]��	I�l��81lׯX5����@s�����,ׯ@|����'?܂.� ���C";���7��b�D��������A���e��6X�<������~'��g[k��ش8�r<������Vz�-O�dhg�����r�30�0Ը�?3H������}�z,��pRDꐈ
�!{S�<^��'N!�ۃ�8� #/�F��F �X桦��Pڋ/�ZZ�iоT���:��`�����ɏTփyz
rr��1����5q#�- �d9���v� �^=C�er$w�_%�ڈ҇ư�1)�,�D��n�~�l�p۬Z���E�"�+e?�̷J F̊����Qں(X�S,���g3kyy��^�_f�ANEe�h�V�^�v��h���}���5L!1��d��I]A�W��^r�* "����G���}�x �]7;�]����b���ؾ�X΁~�� ��g���Y��ׯ�h�J�D�������9���	o�a1�?�����A�o� [��E� �w�c�Q��{?���sm��/�YV������XE -Z��8�@r���l��V�ENN���Q#�|��*���ÂժirsssB�P��,V��Q+�{��\�	���l�qq)��[��9ޟ�/Ԙ��L`i_���;ޏ)dcg�R >�0�z�6� A��P�O~<ow(����U�D�0bJ�ޖ�`jH�����ףȘ�lŞ�+���2~�zlp5���	�Z�0eK�z/0f֝r���|������@�^��߼�]�_�K�H<F��nJ���纒s�P����%(� ;*���5��{����3��i�ͽ�=\����ht��v�F��|�{�,��z�������%������#KK��W%	$D��i����ז��,�s�:�mJ�����c��C��z׏(�<�����#D��Bo�<8����;Z����&�R���֎p.�W>d�KF��t >��zf�*#0��G�T$� l�~y{{d��v�oi ��5Rj���G ������c���aQ.�������(�$�$-��H���>hdYn����sT��l��dm��j'\'i 6�ع�U���ө��7i�L��3/�0����j4Nn�w����.@��0�ȩ����
�a#����˭�Z�r��O�����rG�u���iw)Rk�3,!���a <�)i]q�-�+�������r,͸ދ�g<�Iq+s$C��i4�ߟ�h_#��g��t���!��l���@�R�i�P��K@�Y:�U���Υsa)i���XB��77��}}�_~v��{��\�9gf�����ة����힄��㽒c���<}Za���+u=k^H@ ,����L�ww�u��h�=PkdL
�[5j�����0iTE"1e���CzI��� ��������)�4����;��x��h���fhm]1�Dշ%���i�1�z9kk�4������?%Zɱ��Q�6��g������x�#J��Q]�z���r'E�WLO0?)�w��Y%��2K�,HB��\�4Da0[7[ί$�DGG#7��f�w������_�Խ��b��࿷�3���	0Μ���oP'	;�U��ăΊs��Q;fq
���+����^���n��Ӝ٫歟��d�D�:[˂�X��o�����Y�P����	֮{�zc��U��� z���"�]ޞz|`N'�%��������Kos�z��kKat����q�����#��3�N���1��#ݜ��7�>{�1aL�7n�|>豴 ?��bhC�\YuJ��&9|�����m�zC	:Q��h,�ڧH@D�m'>�)5�#	\�04,�}o�-��������[�33���1s㞫b4�� FDW��}F*-kg��p(��ID����<��-3��V����{�m�Zl�#f���f�}C�v�P]G���K ���\�ǖ���3�+..U)/&	/ہ�$��4D�������\�:�#/e�m��ҷr`d�ʔ%r�F�B#hK�����Y�}�8���;�ش�2��p�Q���������A]� �p�.װ�vGeJ2���i+x�U��SZ��F�jt�Z*ae�׋��`n|o,��S��(%Y�����A$�ra�y(c�Ĕ"����}vM�����#�mm.��(C����	��Ŕ�Ə�$U�uYRJF
�5Z���=�A��w@<��
�`�<)��<ĘGg�C����V����}:[��6PSS�V�T�S���7��"��3�����mqyy�ؤ��ֲva�d�n�՞��!���e;z��ׂ�.:�+�s�I�2���eѴ�
W;�E�o���L�_~��*r,ߙ�	��]I¼�0�f��~�$R�SY�-Z���&�"x<\i�֛��0Mf��&��P�����n�9Z�
�1�@��QQdk�U^^�>�� �d�Z��8�?l���
2���]r��nn��եN
��O��G���a�_��'b��Π{s���8�P9�ta��i�DQ�E���/��y��uy$b�X��8p]eX��|`����\*&�3�ܖ�Q^M�vg,7Y�p��QA�Q�^Ȑ�_ߐ[Q	�{�0L�?$Bُ���ގ1u�ӹ�e:�7b��Ɨ������)흩}��nP�.�'���rd�b+�o'�r�"0��ZaU H��WX���D�����9p��^�^��T[�����HĔ?1�s�j�f�JW��򋺭���%��qI�h%Q���#��M��$��?�^6�j�,Q}U�9��t+Q�����$P1�ۜ;�;�Ő]}?s��O�UV����x�_���bg�m�w�#�s�����J��$���w�.\�r�֦qΛNu����(湥=&n��z����ꨞ�^�����d����Bb�O�^5�����}����{�.a�TV�cي+�����\7�'pڍ_\��N90���?�w�_翍��w&?��*��z=W�~�L�f�{YKS3a�q��'�GG�O��gp߀�/㜆��g���������9���x+�.�4)G�K&�z��b�A���$����x�4���D����7~KK֦ff�)d�$+��۶��{*


��4yUw�ڙ�$ZH�AZk�q�������.�7�#��`i�=:���q�c�]�K��W�T���ފ������,9g�w�g���y�q;��K��cȝ1�kso�؀���U��3e�c:g�f:c1Q�7�w�BF�&����������<�Tq�n���¥<����l6����jQ�B ���hhdo�����>;� l��T�Xd��m���k�hLv�d�s���W[�F�6]�����{Ƕ6sU�@�C�?��F�N�h����kL���&�O`q���{t��k>����U�5I�\��2��-p(C���Z�gנ�����ڜ``��g#��x�@3��UlհU}��Z+��ԂYt�(%��Q-+0Ԙ\Ԛ��V��㫊N���ߌ���xwN�^P�K2�����g4����C�$��5}�PhtAFƃ��׮���[���.�7���z���9���a򡆺�<��(�-o!���gYQi�SA�e\tI��q���� ��!���g�ZG���V��sS(�Ew�Ы�{��2����y���򋋻s��_�1�geee�@����J||�����Q���P���*��Ά��7J B
�C�G*0t�r�tS������ƽ<g�䟓�jM�7u���5z�����X�܊M�t�R�P����"�I����;�%(8Xع�Dw���B���X��+�184��O��*���%b\��A4�L�0�%�t63'a.����8�K%��ƿ���lsF1��(� �R���[�3ZzX�c��Lr����+η��~�9G�e&�Q%k����,a%O������տ�`���\�����}}��������,&�����Y�;��%��߾6�L�5k��5Z^X�W���@��<X��H|Τ[�{� ���J�LXWt鬝��#�Hn��{���/��8h�$	<��<7����͎��3� g(��41�趴��~j��M�2a���E���\�PA��ٮ��$�n�/��&<1}ڴ�#'Ɣ���3�tb�1�7o��<o�f������e
SM���̏~����H�������� Ԕ���1%S(,4�^ef�ۊk��A�/�x�
��q����3�����\�CSZ3��/t�z4��Z?����8��c��sk�NJ��kOGG��YYپ��Έx{A������rOr�'<�9��r�j��ovM�c����F p�!54����.p�&�?;r��?_+��$�䶓SS�=Օo�Y2��4;+��v�``�g�}�ll� ��(`������=qrZ���XQQP����R�yYY#YU���b�g^\Z�hY 3O�ɇ;�yg!�Q|�a1����m6�.9�_'��C
��걸a nL���m~�}�R�/V? $$�oH��@��#�1��������(+K>�P322�-9�|}��D���]�u�\h�^jjju���}��i�Z>�o�P�CdsP�
��|Z***$�.�3��S4�/�̸�I^~���:����ꊒ�}��g/ ��V"��ɞ����t;�KX��3��_=��^��Y�]���pxT�y
�Z�ݫ0���	C!5�������gd�;�q����M��R�r�7�&��ݫd�#Co�"����7�Q�ۍ�ʗDƯ����CWV��Y?O#��u�fkO��W����n��d>R ������Z��,�Ç�̓�
�6Nt,�ā}�:�sF=����e�,�6٪�cj�ι�=�{*f�ך�7�?AP <��V�\���9����X�%s%#�}����W�wy�Dp4觊G]�իtn��&������b���1��-��"V5�&pv��l�P���6�r�� ���9KH�;,��`�=������r��oO��yq��CMU�����6���в���%��2_9J���K����F��~�A a�2��>�I�G��G��s��B��m�V#����bn9�ua�~��&?���$��۱21	E���lk�$d�U�_:
ḣv��x���b���喳�(х.�Uh+�D�hz�o<�b�g � ���yc����[�b�2�O>��a�^__���a<�]�x��a>����|��?��&}����i���R�_7hY�1&��?�@���8^�[]A�x�����X�Evv���Oo�iv�P�Xr_{���K�+���K��Z�a�s�N1�P��;�M�3���v]�r=�}���*����3��u���߀���.]��nh�*	����}x`��]U��{�@�CUE g�e�2.K�� �~��9���4�����X��������,���c�_�����ME�"�#�A�讟S�[q?�{��㖗�V��n7T��2>�**�r,�!vvv^؍755�F311��׏�t����OӸ㔇�@�cp��s�
����*�`�0מ��>����Ci�c����H�d�RF����ş���݋�>�fn�Z�u�Gu��R/:WY���::��:�O��n������^ K�1�D����	R���R�M>޽۶žG�Լf!�er�P	;fEDD���/?��s���XvCJ�J˝�0<���jt,��o�G#2?r�jR�R�!p�_�v�@�4q���{�l�����K�]e����Zʚ�J,�0����>����0�^��1�<�	M?�>>ޛ���(q�m憬����q���w(F�ٹ�m���s],,-��J �� �!bz�D�c!۶�=��p��T�#�Hל�;�L�K�,?�L,&���A��ϟv������
ŝh+]�S+x7�U��2s's�������k�m/�C�iY*����֟�c�{1�$!Y����Yl���0��5��d�og����� �zř����W�"�P�l�ߏ���T.$��7ꗠ4Uh[;�N;����+%�tg��s^�5K/�_���DϞ�;�E��_���`H�h���Uuu�j��x��["�98������L�۠����O�C'�<�x&~�}����S ��g]�:�4CЫ�ߚ�m���+��\�u{]�������Ko(D�'�������1�!�5���TZN=�}��K�/ķ6�r�J�0��7�i�D��ت�=�������e_��7(��$�ZR�W��u���&(<�t|�z��`m�QV��_/�a�d�9#��tɋ�6��Ŷ�"�����iR<Iʌ��A��5�\�bҁ/��� ,��w��m��6����|�`=C	߾)@�K����I�\��J�^�7J��+�\�z�����Fd��S��~��/ᆊ*�~||E
�����3#qq�ٹ��qm)���O����:nW ��ӗ�A�|���{�Sx���Z�t]�
e�<�0�G�{R(��ϜI(��[���jTB�A�!O%3*&f֕Ik	[��l��/(Y�������G1yihj��s�4>���F�����5�ϥ6������Ľ�(������H̥��\ۀ�y�	��^���PJ��:7-��.æ��۰�N�
�P��XCZ�m9.��#�X0��Qm�u�d���D��PS3.��<����A���z�>���W.�JNl��J�Ґ�n��1V�&���^����������LG'���]Z�+@|-�5���FG����.q��L�u����uYwfn�s�e��#���&`~�{�ɢ�I_DDu���m$����EE.��ő�`�U������.k�G�����gDm���R���|§˶t���c~����N�ފ_�\2Ov���u�IPǘ��cs1�a�m��7���ޠ���x�Ժ�H?Ҝ�\=�ma��}�3:.΢ �3N�^\���0)�ۯ��V��Ýw�E�1�n��xxE�������GP�n��:>����)m�6�QM3�2o�b��Ś��o������af!9�����e� p�F���5$.�a�N3����c���<��ɓC��{�%���#�1�p�b��T�a��XD[��,�x��5�Jԏ�t)Z�'�'��ј�������F�PTl,�+�_qHCCc�=+[>4 �Ɏ_�b�Z��������l���|��U/ў����Ӂ61~͙��K*k}? ������|7�1�*RsOP�����m|���5��_�,�ju��8������b�a��Bn���mѨ/��=�6 ��?|�xF��^�.A�j��ՙ�vr^���X4��~u��V��7Ԝ+*�A)\�E�|��'�l�E�u�Z��*�ÿ��|^�,XD��촶�����ڱ�I�Rg��Z}Iy��}Z���\5�+Ub��D��z$ե'��ӡ�P�$��S,z�wV���By�e^�Q�N�U �lF*U���܎w���������p�=ru�˃9�4���ޛ�����8�O(���m��KM^�eJ��{�l9�m��ûq��$�z�$���zRl
��XX���n�+M�>j�v�5չ�׮\�D�5H��� �
-H�e�|��ł5d�B��6�ￂr$������ؖF�%Q����Y�0��d'�՛��N��y�{�k>sQR��1����UwO>E[i=|�N���P��I@�\o}X����7�t���J̕��C2��Z�5C��*'�O�eee"G;S�蹹9A\����!~Y:�Ҩ��ş��r�Q�~'Joi`dgr�υw汹��M������ ��?���	 �kB�6Xiܷu��a���3OOo�1�uŀKoc��w?;ڜ�i��������M>\�~��0�B�P	.��`�Ք�[,��4�@�i�(�kdh�(u�}�q���ӽ7��i��G\��C� �T}�U�][�h��4���QQ��ͭ�e�]%��k�C2�v�S�4׭!+x&�S\�@�s��ԯ�A5e�>�������Ju Q6C¢�K�»C �@Ã��x��&�&F��^�OtE�}��x�����=��?�M[厦MOf��וּ ���ck<�ا`��PYZZB��Z9e{��cwfh=G�`�����k/��,}t�?π��� ��]'���i2��.�j+���e��<�l�r1���n�Б6n�Ⱦdx�t�xҵ�BO��?�����o��\\�Um��E�/)�^�V�
XR�'GGF{./WTٍ���-y{�n1ݝg/���h֧��cvv�Nq���kp�^�cv��X�'�� �y�`�}?�V�b;k���Z':���Z�'b7�٧b�e���a�Ϊ��Μc#�����+*B�ٔt~��0�hm���B�-����CV�5ؒ���i��|�m��3{%�#�|P~P�~Go�~DDD�γ>�]3��c�z�����Ei��i#��Iė�������/č9xO'�E2����ѝb��a.�X����/M��=�;�e%5(m,�r�T�Bڧ�����܍5:8��GGG��؁YX��w��v����H���
 q���:�^�)b���,z�n�}kԚZ�ۣ����*��*�����x��nǳd6�,SJF^�j̎c|k�*[�����������O��T�(&�w���2�``(��w"lhU�E��#�ڰ9�Gt�t��g��-f�����B�m�b���&[;�X�G��mm�3^�$49 ~��C^}2#�h�o~u����әw��D�h���� `�5���>��%����W�o��eG�� g߾}�1�꼍u�$FEeA-F��!���&��< ��XCBU#.>�Z��j������p.շ��� "��>�)&�ﻏ6b���-�W�А!j���<�z�4XKĘG��RY���p�t�JS�8g�Ϟ%�d\�
�l+*�?�L������jx՟�u3k���ׅ��L�bao7��AC�Ǘ����;,d򑉷�`��}�.����@a$�+�&�@i��k�4)6�x���6�]p��U� £s�4Ź_�+����BF��!��&`7b8%�^;� �Qi�y%%���P�h`	�Y~^�c����8q�=���|9eeD�
��+�::9�簾'����!�D��Oz���,%a�ElA���jq7�go�߈�;������
��Z�R'^�����W�^�D�`G���?�H�X�/�k���,T�'���F��R�P���0o3�ۦCW}�.~(e=��D��4}��y~ԩ�%9X�4wuy���*���K/8�k�S;�M��@4z�#~|f$� xZ�xN�-�F~�n�P�S���f�ʭ�K�_%�b�Y�ؘ�8�acc���"5x;�?i��DI�(�ߌ�,9O�)gp��Q�7ܦ��m������;b�o!!iK��m��f��8`�n4���97oy���[p�n�~�O��O�/��*��}T~����e����O��&��X	1��r�~��g*�]P'��4�Q�U�_���u�6�9������z���щV�h2�Y ��A�<��_����ׯ_��g?]�V��Nv�Kv[���D��S�=��ڭ�~��A��9o��=ū��/�����C�v:�$�V��n\�u_��3p��
F�#���;-����Qv}��2ڼ�ή�E������k+����?o@Y+�B{w�2Z��po�S_&�����s���މ����vq]]���E�z�,o��a���RDD�%싩P(�h�^��#�����~��&�^�vc��~�X$'$���������L��*���J�zw��L05X�qo�b����F@�����R2�m̽}kp�o}�h	Bϟ/5<T����_m2�Y���i�ƽ�fл�6��\>��4�Е$�V�t���}C@@Ӹ-�Xt��eB������t�������`�[�5������X�Z:��.�#Z!%��!*��j(e��_��s|�4E,���̓����u�X�������'�,��P`��G�5�q]��v�p���h��Pih'@�L)�UUU���
��1@g��zr�k�	cl���c�Pgp<�9$EK��89ݰ.� p�<�JnPpp82G&�^d.ɉ�uI;;7W�cU�L,�{T����^�-~X��vZ�;*�m�c`j���X������*@������d��~�,1��旃:��G��@kUiїaV��M��E�xڪ^.~�������zΰ@�?5-�~~؍�S5~/�r��N�6@�d%��@�cq�E6��h�9+��~
���2���៉B��1<�T�#괪*��5�U�99����~�hF�8��Eѥ�����eJ�����,Y��(��^�}� ��nb@ðid��,3k���|3��_*�덙>�n:ևz7�%������5��E��~bjj꧝�PL�i5ߛ^�����G4A���*�F�.AAA�:�]�~ �#��+IJJ�:�$���q��ˣ�v	�`[ۏ �.\�k����рF�v��p��߯�{���-y}�����atR�����#��W�5�l�w�#=O)H}2D��g�n���&]L,�0_��
/�NH�䐵��T2���<�}t��O]�����;Tl��{��1e��a�:�{&V��|E�Tn�� ���#����=X�8X���2-���Й�2���U�����J�l�7�������5����j\�Z9�%��Yf ��ZC�hML����iS3��'��)B.-�_�����r
ҍ�</~ �q��g����B$w���&�����S��"�҆��8����;���*�P`D�8\�뱵D5�<�]��U��,���???�W����$�w�y�l	P��ր�Ϯ)�)",��·ՇY"��#_<	s짠͕��@/g9H���4��M$�ώ���w*{��� �>�q۱E
����c�|9p�,˨G�3;D���sY��W:+�-����UZt���L#����׹D����Ÿ��~+�S�ɾ[�wuw̯��y(?�z�©`a��q���{��$���J�A���� z��(ʶ��çO�}7�,!�Aع�~%���D�6����oC�k�B�[�h�������|�j�#R�H�D�|��!���ˌ9��\t��ِ��p��=ܿdܰ��1�72��O����"W��)%��l�5�o4�����{�9��
�Xϰ���H����-�=}�w�}�ۗ/�y4$8o�t�٥H�:�vA��)B���޶{^�	���|�AW/nDr��mQK����i,� ��)�#��i�~��ut�7����G`%��+�ak�P��y��W/9洴�pP��h����t�7��3W����%�ħStU�թф�7���*�K�kM�kb}���\�E��!�(���� ���Y��U�(dS���Ä�UZ2�s��s����[�2PH��M�vK��JD��(��ɟ;��J�kW�C�~*���1ş��EP���-�X�Y�)�C(Q�*���S����jjhd���>�`_��4ڏr|��[�=�+f�� ��������||�p����6\�j���lؤ·}���_��U+��v�mX$f頓��t�K�/S���<A{�0N#����yt&�wA�рqcw誳���r7O�v/i*6 v%~Ԙr7���
l`.���eg'�'Y�w��T��@c�W�b]��|=�>���: +G�(�|�r�3d#Y,���7$|7QP�:�����To��Xnt���q1
���1�BN��:�4��c����N��c��!�N;1��+�kK�@S�x�	����1��C�{Q����х��TŬ�<����Dj;��0�`������	�>�l�>ɖE���ܾgn;����bȟ$��>@���_��h&��J/�k���ߩ����-�E�zaº~�)����1v^�Bå��ah.��u�J�
�������(6��ł�Oo���Qq�	l��[K}@睻p�Fu��e����'a�ӈ����x�'����q�r���E�8"l�z��GJ1w�?RQGw�*���!�ZVld>�2���ph�����W�sJD����� $��"J�JZ��$\�r��w�U�e�&+Z��~��O����'�s�� ���(O���..��VL�kih�IH2xo|ߛg����ai���=O�i���`Wd�/�ǆ�KD�lOߍ�8~�4���5��O(���~��&WʘC)�{B��v�a��'ڥ@;3�C�O��w�}L�;:9o��31⩶fA�!��Q
�2K�.|�B�2Ԋ� Iu�Q�w�b�3w(7��i��R�g��ְ4S_�ؘ�iQ�P��5r�Q�^Hqڷ�sfD[��v�G1��<����m5�Q4�$!h�rp��hTu��Ǌ����*�?��M��x~q��l�g�Ib�?Eبs{���{l���t���ԛFC�@�K~������`Iw�<=DZ��|�^�������0
�V����E\�jjj̖��7o�a�j,X!cjk�8���E1>PR���t�$Z���w�Ξ���	XO
W�C�����-���%��Wd����m�^����Uz�4�hE�̩I������f��j �B�딠�7��x���#m=�ͦ�k�����!�]
����	�u$og<��Żt����G��b�����'���T����|{�3�e5����B�T�e]�8v4[���~�����"k�Ey�v5��z�i�x9����zš�JG�Jp�V6h�Z.l�L�3-T%����@�طT�������$oW���>UŊ+��-�*����܂��h�͛T9Y�+��Y��t,ߙ�'������|uF��v�m������rB�@�ʊ��dfa���RQ�1��2��"�������g^` ,q��$�]���������eeT�Р�p-�5A�i4
5��e��Z��o�3�j�J'}� Lɲk$�>HQQ=�����+k2�����V�^���D~�f'�cf�H�[�N���m�y��L���j�ԻV�E�G2-nw�n�`M���M���E�d���
�(�dLц�'���J.���6t�^��c�VЩ�J��4y[A���6^������I��z�$�W���`(ȫJ�R��^���B���F��c�ys�o��Jg?F*��0��?�~��N��C����w���F���F�N�ɢUNsJ��7ђ��&'�_�v���dgԏ�7��f��O0��u/:Oayй�����G�Mv|w��Vl4y���]ZY3�`1����{���u�2�[C����t�����%���<�=�OD�0-���Z��n���&m�m��"y?�G��O�xގ��b�7z�S�k��'>����ȝ;SL]���n��t�����1�5������f�+�FX��^���q��ѧ�0A�q݁X��p���`���*ѬH%1��f���R��y@�a��ٗي��欟��o�x�&�Œ���k�iД���0�@�P)/�qt:�4��!��ɯ?����-g��!<�C��Ŭi�#}�3g�P�r����*{��%��1�9y#ݷ<�s���C:"��$��Iņ<s�DWZ�w�\6�7j�Q�E�&M�5\"_O��Ú�dC���_����:�܇�[+�S��]�Ll/�$��39njj�%�7}���K�Po��__�<��2���{���}X�+k���n���*Ņ�p7���bu��M�mV.��,����u/{�㥊�B�ѓ#2e�
Lp]�_�)��>�k�*��縇�8nc�<Ǥ�n7�>����H� 5��mf�f�]S���=�>dc�����Wm��
��#G�d��ͷ]�PM�i�3+�N�O��W��8�Ǟ�#���=�~O�[ߟ_�<j]�=�z�����-�Dad�VƊo�W�l^�g�?�ua/��(_�hƳ�Y��Wb�FNn,���m����Fj��0�x��虧/W�xļR�qC����h��������8l�8�T������c^%I��s��c������.��K�q���ϫ���+A>�="���$�%�r���]�1߲��)�L����1���ҭ�Q�y^(hb����r��q_�q�|J��b��W\{Q�(>~�"�:܇2�.y%l)��,*_�[	<��AH�����ҕh��������Xw�<Y\�KI��#���=�9��g�V�_�y	Z+��e������Lr�'G�Ep�y�-^F)֫]ۇ��jY���va�ha�8���5t�����94��.|Ѿjfa�nCl1��8T�6 ��P�L�k�:n˭PqL)ds�ՐT�0V�2t~Hǉ��0mwu�S^z�|wF+֢���K���3T�z�D�1�%;<���$��pM��D��(�UFX�-G{�b�V���%�7���j�bX0�`Qn�l@����i�24�(�*���W�|�A�b�v��˫v���������qNξ�P���Vt�������]km]�n��Q�bIM���s{Ɓ�CA�6��B�G��Ӑ�����Wi�N�q&'��S~�s�2��w6��3��N؝6�+Z�:���oc��E-��Z)���4�E@�
�0Vߪ�5�Z�-�S���
=x;l����K[ ^�r���{��.qD���D��k��X��uU�3�bH5A tޕ7�w��¦#pʫW-�7�h���L�=�w`E�^�b���md*r��l���\��ә�[�cm��ϴ;_���eR���B K�+������%�]��+Ҟ����(Ĥ����s� ϞIn���c�����1�
�acm���?n��o0b��<*�g�ض��'����XyV+e^��9�|G���x+,�nP�S9��+0��?��fߝ�Yy9�����^A��v���������,��_����X?5�� Otn���It�H`K��s��Z�Qd)�J�1l-�vy�d�
soi_d`(�մ���u32�<��_��n���'9Ēn���{L�&Y� � 6����4,)�4��۲6`LP P�%ߞ��ʦ���,��%���q��T���3���/1�3��g.�s���5N�9�Ű�?���v��L�H�6N�ϭ����@;􍋏��W���Ћ~�x(D=ո��.{d�z�tYL�rC���G&�j�,ug
�0��q�����
־�;��<#;�X�V�D[�[��[46o<94��Y4�f���l@�H;��p���nrd{�c���l		Ef�#Op�GVsD���.WE����.�t�������Q��S�-��|_It#RE�#�n��bI��6�|�Yv6r�&�O5�Rh�i3��c{=$o�t��r7��.�w������Y��D7��l���WZ��E�.��� u�{�]̿%��q5]�Џ1N��$+9�f��?|�Y�'7DN2�gK>kXX����2V�q��/:ܜv-h��Kg���H1<�>A��Õ�1R�O���˚`�Yk<ᝦ|��\z���LA��x?r"��T�7��y2s�У��T�h?��EW�[��/ghX��!�閌��5J"��A�!�$#]:�r�0R+�bٻEt-��p�59F�}�Ϗ��������cco>k��R<O(,�o���ˑ(�X����l��.��>r̻d�@��i[%����)f��s���m���^n��j1��u���B�9Z����5u}��^��@fG��'�_�:u(2<�_w����G|�р�Z���w�`�1�#��j��b���əZ��C��Ag��O& �����p<���D@7j�)Ж5�r>��wf�ʵ>%	�b�jz��y�>�7e�c�@V��!��y|Vw�$0?�b���-��=�mbp���+r&?&����D���ʿ�X_T�;�!݈͜�U^A[/�W�����,Y�k��=ٮҌ�IYwc�v(��a�\���+
hFTi�)�;a4�X����O�Q�����"��ET�2�%��d�a� ���֪����r=�N�_
�3�_>�F��Mq������wy�ҡ�'�dBIӆ\��U��
���?q���u�R�5i��x�"�V�H+�
p����/�5�G�x�[L8���W����混\ʖC*�3�(�*�C�ve2�������뻜��,�tJ�3kWG��m�"��!�K����Y��1���9qSU��L��-��Is�1�K��~��]��p�Q&a��gБ�~��w�����)���W�J@71�x;� �RK�{rXѣ/��."F"�V�����GZ6f}����qK�����o|�:��ϼ�X��-��WۂzpE�w(����Ɣ��V�I��J�v�cg�M�ݎ���_<�C ��N��|ϋW!�[+�_X�+�����$!P�Y��%Ӄ�m���@Qek9u�z8>�'=|�BVK�c`c��������T?S�b	�������J?���D��G�qBK�n��gm�v~�f�g	"OT���5��g���v����d�DWf�f��F��d��8�_��|�r��L�;�B⁝_�WB�{��R��9��3�����~���ׅ��ۍ��,�yϫ�֣8�e�Ѣ�|����]d�n���_J��Ed�/���2���(��7K��e�BQ�W�A+�K�(�b�n��G�Y��)����������6��|E��
m�����|BJ#�.Y�௜������:{2���u'����t����74|E�GBM��v�wS�,}��yS�����m���QF
*R-|�?�SكS��۫��AĬ�7�A��˝��$xٲp����X�0��6D��y&K;��T�p��:�r7h=)Tv�?^�%��3˷Ž
JK�	���E�;u4wK\��d|�B���|���$9�-��{��ذ�g����Wc�#�ԇ���\;��y6?	����h���>�c���#�OJ�C��|9��;_IV�l�m��ܟ��S<p�c�ںz���G�5��p��A+���Zp:��o/ߙ���e�H�Դԙ�����n)"�i咯J��D����)��~~�W����8��.Q����0�Eo�׏=et�κ���q,$+�)v����ce�J9��/5����V.�0����wqR��%}�[NHɲM�_˾/&�ޢ�L<�z���G&
��Sg~9���P��X�H�K����M�R�GЕ�{�[|,^�obi@J���]{��t.�h|;2��~�F�9tnsIRuk�w5�	"���c���K�Ƚ*��{�}���uRM��CcxB~&}mJ{֔��'pS�z�b���l�O�Xa�Z��vp�纻l��m;���K�R�֠�h�_Ϝ+1���W������-~G'V}��Y��b�~/1���,�Gv�f��5��$�{�ə^�s��5�µ�b��G��+��A����D�R�W����=���������ݵ=�;S�/K��DpmM���7^�:���{~J��9 ���O�4�*����W�\փ7����SӹR�Ɂ&XcP@���UW6�� q-z�#��=?0���[Ra&?s��3Ȋ�4�����X�G�$���>�"�;Z�����8�\�h,WGWؔ�$}��mΑиy� �P�5n��]#;�I�L٫��=Zym/yc���h�ъ����_��A��W��Yu��/�uÔB�ʷHgX}�kE����,��v�fk,m����UʡnB���֭�}�=b\g2���!Js+H�vL;¤O��ZK�-��_#��g�?�DڏPS��D��<�>f���g��K��K����%�&�܎������2cj[��F���mأ[ }̢�DE8�>��/��2����K�o��;5ȅ��-/���֞\Gx��P)i��;�;��Bm��#Oz��<_&�^:c��#$�N�KZ��T�u%�n��^7��4�[Ib/�0J�?lg���YY�?��un%Z�"zN�y�*���gBFGy �x�8���y(�c�ԭ{]������$Ez���,-��2uO����Ԗ����z������ͭ�2�|f.�!�0��C�-�ŭ�OՖy7���Y�m	�47���s��~KL7J�xJmw|\��N=�������(��}��P� σ7;�^43*�j�Z�EHфzDXj�����h�\� ����hH`d�"�L�}'GIS1�
��~��+U'<�vz���K��h��?Sp��O;ig�B�&{�e�z"%5����b,T�!eny�B��n'�F�x�*�Dq�����Y�E� f�6�õ9>7c��8�
�7�IODUu�����x�^,�I�N�T����Sa0��E̛&��˩!�0�'T"��/��|�����2m�?SJ�z��XL̵4b�޶ݡ0�Z?�m�;!c|��eW����&۸*�t�|oo���c� w}�~�8����<��b�Ei�C܄IO�Dߔ�_w3����<�}�~� �L��3�qY+���TP]*?a��~�>S�냳)�A;��$�^H�v��>/�ft�bU �-��iWٽu��* ~GjRs�X����Ğ`�Ocv&�F|�N픵��ut_Hq���7���7MFoG��#���7�=��)F�}r�s�3+������Q����qU՗(���V��Π�DS�V��
��w�ė2(KQ��BY�6�e@�z�h`ۖ�����q(}����� �r�އGQ9"�
�������0� "�C"�C�
JJ��P�=��HK�Н�~P����?��\Gq�yv�u��ޱ���@w�O�0��!e�դ�x)�� �%����~G�m+SֿcD�)ǒVZvԔ�*t����Ė��h��%�z�\�gp�α�������L?©�5}~��~����Ǟ�f�)�L03aݗ-�n�':��"�"$����n���U��:y�5\��a<ܳ&�y=���t�c�ܮ��KJ)B�
l}����ģ��k�D{{s�h�?>��ͧN�h����/e�0�t�Wa�󔨟���,�,LU��`���"5�Wq��m5��v�]���Kh���r%U3�Т��6ZQ���x5�Ek��Q�<3S�e�\�A<���n*3�	�t	�t${N^)Z����K9[髠[|���SeN��+�N9�&��f�Cts������O��;r���z��pFL'55GY_y|���������2%e��ק$��33Un<]n�	{"%�$�x䢭�x�sr����²(q䬯���F�ECfD�wh�W��F��e+��馧���mp4�~X���2(��;��n��'���?���y黓�{�����9*ˏ���D�DD�?��~=y���ۮ�R7N�|�#���_[g�˧�t�>�m$'�h�u�*G�F��tZ�!*a}�.����N��sŀgޣ��s_%}|�t�Xӿ�ݩ��Ԓ}���(��b�#���k�b-lY���j]���{-��iO�$���'6���-��������ȕ7k�9��ST�6o�#^}�67�֪��	�QU�JZKE�N^̃�X��앖י$a>P`ZXT�=��E�!$*
��"��u[okk{�
�����O��|�Z﹞t��d_�9���������ʗ�d�	d�� O�RSM���<Gax��X��l���� ������)6�?!�����h�η3;�͆�<�g��8V��qV�*��n���R�^����OO�~�N�G���4識�	�����]p@C�4��>W�`���;g;'>�ꙑ�J�!RIv�rJ_�5߇,^��-�KEdk�ol��Ő�_na7��2?�w��"��gG1%%%��8�F���S+���ȣ��67��糐,Yʆ偗����#��E۪�;�g�T�
���4t]�jڵU'�Q^�T:y�Ŏ<�nw�ל��k1��%�1GA�=s��r|}O?n��C�����������E:H��RƊ9�EO|=龿�;^�:�o3����xW�,�\wg����t*��cU�!����r�;ꍯM1L�йp�d�X��ϞV��v}p�������$��3.r�,&�h�숖�ꋲ-��7��z_m2�1�p�e]#�y��Žm��P���[�����ѿ����H�n�@���[����U̐٬��2����M����~��]g��L��z�;��c�xZ�|��Bx���{����m�$F8'��"�a/���no���ew���C�����@��aə�H�=�����{O�vT:�dcg�K�i�$��z��qKJu��Q���)�@b�С�T��B�p�h%v��:e^o�zΛ�J��ի�g������99�����i5�����g3126�x���{8_p��8�:LG�^:�ly��ezBpo����z��Tf�2_� �}�rm�D~̩nS.��㣍�X�C��P�1��-Z�n�g��v�x��:.�|�bΔS��fOr/���SU�q�	�癤�Aq��2��j;�w֣���6:kI�3��1�8����ڶ0(bQ��4?_�j������B�?�GG7�bg����pw�t^"nV�1Gm�v6����i��W-p�:����UG��l�߫x/XK%����|�;}��Ā��iB��FP
I%�J�j��K����o��HZ���9�N��s�MJ�oX�'��^N%��52����ٟ>]y��5��ٳg�deU���P�J��e*1�󽳝I� �����}%�膙z��N3nͩ�vF1k�YE1��dnH�e���R��T�z��~�؁�����VlG��D����:���X��[�x���tFW�L�s�q�b��MwC���܂$��c=����W��������xQMc=_mix�:+.-6�m�߽���|_�f�-�Vz)))��ϒ.s�ƨN�(?�f��$����l��G�s.���p*dp������߿:r)|���Q�]"(4WUQ!ϭ<�0"S��.de9�O��up��V�$i~�H��xW�QL�~7BG�Y/���Տ����j?z�X+F~�����+��\c�'A9�A-�����5��pB�^�3[��p!\��R0$�|VVpe��
���)*OM_i�2W����8�&$̬˲xn��z�j���q-&뤊㐰�.v��k݈����{̓���;�B���;�~f�U���.]�R������⒒k�q.�S	���XM��@C�]dӆSf�ˉ���Z	OxE2�ߗQԽ:���x6��5\z[h'�j4_b{�.
�O��ʦBBXs�:+��>g��V�Z�ІN���H����zO��E  �
W�"̨!�I[�g�;}��1���������&(6�����t����Ԫֱ6�����i�Si��L|��U�9�
�z�06x�����!�e-�������#�l7͠��5`'�\���5�{Xoc��;N���W�i�SSщ�5�#I�p�_�Dn]��''�=/}Æ'���Q���M�X����r��D M�q)��,���������$���h��̿��+)(���w;��I�5G>IUԷ�*hI�_�G�j�:��MR:NTy |���f{�q���M��WMM��[_����<�<łh��ݪ4Bn��e�u>����	.]xC##3vv����H];�#+���`AAI���@GG�x��C������V��s*UP�II���Ϧ�)�S��[��54"���B����з�" �@׬e#�z\���Cm�*��߼�E�
@�"����"5es�g�!�zg�ݴI��Qzy�L�rv��͛*e`�NN�5��t&5X�k��̏�/��(��#�a�T:�a��2F#��V'����}������ԉ~� �ڝV��\a�S�� ��7��4���֚�(}��e�g~�JKKsVB���F*J�5\\\
����r��[B�{i�h�GN{ss���`�^�����(��껲�&�q���Ї''0ؙ�i(������Z�,���	n���8�,�|�ljr�\J����6�(����lj'�<|v������8���g�1ek����w��^h;��?>�EşS��aa��H]'H����g�J
��mJ�|�F)x��\�\s�=�T��"��>&�yn��s�����^=*�?�IFKkonkˮ�#�l-�|	�ϢUt*S�ߴ�N��zff���`�i��Y�MLL�i�E�Z����1}oK8�>_�3�:��g-�o2���µ�YK��,@�m���U'��C!���Ly�X�)H*.�P:�^���X͛�����C��tez�� ���.S���F�Ħ7)-�Om`�,�iM�I�c��d�l/e�T��G���$֟�n��7o
a�ast��IϞ�e솲_Co�p��qy@�ϫ���� Mpʔ�٥[���Yw�@̇t~P�����4E*~�����N�/{�+9�))��};�P�`0�DK'.0ޕ�.���q��)ڙ��Sf?�>Xמ�t�̃Q��l��Š�)@���m��5����U��Q��L��?B�.��r��Ȥ�.��\�%[sNŭ���=J&���
*z.pgCqqqӃ�U*n��v	t���s|�3�ɝ�d?�'�蘘�eW�I鸭�A�.
���`�fS�����D(��Jj�yp��6�?"]�e+���p=	�X�'�ɰ�)�٩|e<+y+�5��l ���m�U��[i\��V�DIu{���b�'��J��m�5���T����Л�q����έ�������>�G����6���8�h��"X���gɠ�]�Q<�>��٫���[=��{x]�P9֊Q�n�'�D�`sX��]�#��OS�2� &���	]	;i+q�L�N�Y�0�I�-8s{�f%�;�l-�gt=4d��:�����n#␕=��L�S�-_��݋�}��Ĕ;0�=��jA�MN}C�9U�#�th�(cy0�$,�}���eK`aӅdq ���d�B����_K��k;B�ef�+74)g=�S�H0W^�)����PϠs���,��W�AF�;f?{���2J@���r��{���g���od������ȶ����Bw�N��u��-��<���X6NH:�Ƣu����㊓*�cI,�I��F$+�_���L]�vH��˚w������R�G�JO��(�D;G' ���B�#t+L����ǏD$$��6_@�X;G���ܬ�CQ�y��F)���<���L��6g�1ܘ]-��&�_��`,�z�;V3\�Np]*� l|����I	 7M*2==�e.9���T�],����`�u=������D�=��w���:���R���u�Jlly�E>h?��&��o����y'�����X�Q^��7�v�^rY����xql�k���� ���QRA!�>�!�4�=�!(

��B�$+�סZR����e�*�k�
�������y[[����@�dC �2~�h_����	����e�&��P.l�h^ņ@���ii�j9���/Y�v��a�L@�2�����g-∁
	A��~�e������Nl>r{��)4bU<����Y���-͈&��a����#��]'�PS4�j�f�o�U�>��o��e�ͩ|5"!a��8���w��SOp�Ƃu߆BhF.��~��G���;Tj�������OxC��I~^^Hh�q��h>�V��ݦ��ϣ�Q�۷Š��s����G�gA(�L9���}��0e>�t� J�W<�TW���f���������@)�#��à��#�TPQ	i�����k���4���$��c�<��y�����H�e�QU;7����{����4h&��8�o���������z$0��F���~,�3�|>Z�?�c�w��Mff�s��uҺ�(\\�|0�$���X�X4]
������'�.�N뾡hYw�ﰥ����wƵBJv�����%^{i��O�����D���;�?~�o�v�A�J�a���m[�0�����n�.w��>�<��./����Yٗ�5�ώ��*֒��	U�xEH�t<�oM�[E����eF̹��
�M:m�$�nR3g��������9ם�O2�v�@��I�y���l�_��'#�A��&��A9j>E˺��K#�aoߺ7C5ej�;��?��V�4:������o�Q��"z�||@�� �`&��:�����	a�}��B<p�^������N��ged�EEEe����8w&<�O7��f;b���� %]Lc���puv�m�uo�(P�#�디�������c��^t��ӭ\Og:ߗ�WP8<UhgkUs�\�9�(D����/pT�����歳���Z��rX�����Ǩ�E~�����Jy���n�e�6�9���,x>V�$������/ĭ.��(_��X��%��p�[m�.�U�����c���ɐ^EFj�H�9�,�������//���:��(�0i%%%R჎���V%/l])�]�»ahr�f��f�z���A����2s �333+��������4⺜�(� � %������0l����C��T�n�Ny���0=��(�vg.���j/n����z�g�O�r��JHH�W�k�҅��bE+BG^
�ꯡn)R�6�O`���J*�:	�l�C)� ���>�~Ip�x�oݥ��f*�����N_�#������UH����d+]69b�7{�;�\����i�����B��j� ��I��K]3-��_���a�m="н��XHt����٫�9(��y�c"��r����P�'vQ���O�7�g~c��:W� ���Q��&�<�lh���3��@�#cG������O]�<,ii+|�������ի�1.w\�n�"(��ǹ%��ޝ
�]�^=�� ��͆�H8;;;�� P3��E�����Rn�̠5�;&���'�_�*:�}���~��Ya𘘒2�>F�?zA�x������(Y7\��}A kX��Y$4����3va��P��3�����D?ck�>_������, �O���������l&���lb�����6�	��?���'$$t�z��7��B�I�7����?g�`�v��ω���'���+�ڿL�O��w<z��UlUu�����&�ݻ ��!uEP��!�����"���KG��	@AG��v���!��v`�@W�����K ��=555��V��z}7��p�&�����ng���;�2�IL�խ��6٩�t�?�"6��>�e�)�\���kޯ�W��'����^I��~��Z%m�L,�5K3������W���x���Gh`7 �e �)��莾2#Ϊcp���fLh(�	+����d�p����֜��H%�N�y1@i��OC���\����{(d?����o߾�Jw\�p���`bb�����+J�?~�C�5E&^��]P��0�Gy-NDU:�g���ݲ�
����U�T$%�]fվ�������2�R���D��ds��e���A��o?�@��C������Sh��Flq�;���Y*��ۂ���VW� �I����4cFc�{��A��ցG��_�N4L�:��àZ�ȏ���Y�'r�h����\s4�V��?O���J�ҧ���> B*��c�A{O��H�Ha�*��T� +A��ai��(҇q2�͛�j"���|�N�2v��Ȩo�
4N��v�0��}�t��v���<M��o��u�_��G�c܎0�-�2C�Wy�gf����C?e��)gBȞ���峀ׅ&���E�9n@s�|]|λ�A��Y+��޽���-Y��+�������R�Ӝ�Ν��
�Ќ��؁��1{xV��!Tn/>�w��ֆ�
x���E��ԗM�m*�?�0n[
�2ƕ����H�D��Ѥd�9���c�h�Z/Vd+kQK]���L.��5�P��}�9pô�.�I��N��{�bon/��K���R�(fm����en5��!M���Y��$���PE�]�!�}�����:g2�455��@:�A��~�>H}Wl��T���ru�������B�	�`��:V��G|jS��c�@s=0�mk�q��2����Vk-bz}�0�o��$pQ�æe�+d.0/��w�Jcݓ$�嵜;!�ԙ]v��PQ��,�p�A�"��%iY��ǼO���:ϫ���?�o���?�N�Z����AiD:�cR�?}��9�������	�)d<6�4b6	��`��);۱A�>�^�ΔT_o�/PE����Ў�,%�g��N;�_�-<���k�(=g��4�Y�*Ğ?��͛N�ԄQ��{��/�J�&���ګ�?�F��-Gӿ�W�ɮ�ʟ�t�`m@����F�������2�33�����-��Ш(s8t��Kr�0�袬Ũ�H38��FZ; �Ƞ �	#�"S`8�w{�Z��s_$���`�J��)����G�Y������^a��S���RJJj����-'�δ��I�����3��MEG_��(wX̨���u�ɝ�1��(S����|�fN
�����MvҊ	�گ���58�i�<l���>�����i�9��/ t���c��|�r�s��K�!��d|jk�_� �g9��.����:;`N�TGc>�2��aa�	�ouuP`J��e�L��O�s������ϼ�g�8�v���.Jq��w�u���#��I����󞧷����Yj7C%�&y�I@�XRRו,��o�,UE�7�����޽{?]U���S�y�ڀv�_�D���c}���YYFF)�l�������y��h�k�N+�k��U��,���Z��Q����J�����+˥'a^����#%�v�Z0��B�.��B��1��3� (��ǁlLL]�g�i9�d@�����:��2��׀���X�q���M�$s�7���nb��T�%e�Mt`�d�9|0���8��<�hg��o6U��3wbJ_#B ~�Lo��a�1L�Z��B�_�f�&�G�4VH������[��������x�v�ܷ4b���9c �̫�o���՜c�\�ǹ���� UJV6k�z*ݝ;P}� �k�Sd{�$H)()��h<S'��0�m��N^T1��2M�}���cL�n�U̜��'I0 �CK�s�y�$�
~���t[V�}��"q�g`��(�щ�V��������%�t�C���B^���{#|w�e���p�M\/*l����)���£�1Vesw���`MH$5Km�M���y�.!�͞�7�0h	��ߺ����W�L�r���s�n�J������˓q�++�ec��R�vXǈ�?_��V*Э/��h���k������j2��=�Q�툶���B�O������m��^��k-y|1,�-E�QӼ��n�"�ksp�l%v�5q�Ń?[�T			PY[T3K�N�R������M2���-��>����l�K]	�UK�@e�(+>^dnn.e��Y�gI��^'0�J<ʬ�3�oM-2 0g���}������m;��)k�h���i�[�k�������kx�Mb��с�����d#�^3�6ו5T��=��H��5
�b5��+�{��;}�˯��֋���S�(����1Y?��UTټ�R�I�D�YX��0<q�q�\�n�|eS�Y��M?��^��0=<�E�,H4�bI��Yu�v���YF��(��r��o�/�(�Y:�=.�+d\�(Զ��.��X��C��^��Ք�>�9h�2ٮk���ߖa[�W�U�+��Qop��U�VT-s�2e��B�r�՜�=���&������n�O�Q{l��r��c+W��e�D.���z#�Z e�܈<D�
��J��2�A˾����-dgX�Un�:�3.��ܮ�t��!X�&�$>��<2b>��'`���ޘ�^r��$��+	Ə���ѣ���i4�,x�8%�))�1���n���P��G�?r�^�V�A_�iǂ���;�5�%lv����R���i��A�L���vV����xI��{��ݻ����-�5o|% e�Us�E'��>h�3�<���k�������w���|vnm�<QPN�B@Z�0y�?�
������5_��G/�t�@�DBe���0�{�q��M��xh1���9U$����6Oq]*mXUlH��i�}�a&;�@��#&o�8ם:o��w<��я߬��U�y�6UZ���=t��+����g�l[����I�2��u��3��}M��T��*�g�[�*�RD��i��V%cg�R-��/��z�QY���wA��}���Ơeh���5>%�E1��3m1R��h�> X��q�EP*d�V �!�n(�;�[���˗��8&;��^t��;�NP�)�� @4����񵚝�~��2
@���DF
��[��aa�tڛ�����T�<e?���\�)�ں"�&~��T�faׇ�bP�%&!��e;���B�;��A�YP�N`?B3��C��M��9T�����9X��
���hTSQ	�8PI���;О1�������m���@�4дR22*��/�z� �7��>�:�B�6���3qK��wZ�\��R,U��ٗkjB;�*����ʵ��j���
L�d�,xL/�SYo�o���E���^$���M��RoL��!o�R�6"̫_�>Ѹ����R���9��wo�v�0r�����(D"ev֤ФST��~���6t�locζ4Áy<Z*�b��J����Y��hO�he�A�29�22=��
�B#��CJ{8�\�l��p��T9}f�p�ט�Sx��;72�>��i�|��l`��鿦�����%��aHT:o(���Bu��kNe�cY19�22-9��{1�>�p�'t�ǘѪ7?/4:~�Lù���jO�Y�u� >��4A�p^���;:H�U,0鼥�4�*`���t)�P5�a�(s�b��YfT��P��٤�=績LN��25]G*�G�S�b2F؎�0*����_,���v�r|�����L��] ;,�D�<��/�y��k�9�
��q��/�9�\��=	b� ���K�Y�E��04Bn�kx���?F���O(,]p=��ۇ��.N�6
�*.2Q9��ʑ��T �A�.�p������=���U�g�� �P���k���C �鹹�O�c��	Pt�v^���NVU݁��f_c0=�����!L�)ɦ �4��	iU �&"�;��J@q&Lmu������R;�[K��(���S���`d��
 �z������a|��}��M�Ѝr9dԮ�E7&�r�#oc�bX���fYW�>�RE��x{cg"p.D�^DM��qM��E _�XF��["8Q��=&1MN����� @����o�/��A��=\��@� ;�K5�o�L��E_rTL*�#�o��T�*�q�[�`0�P:h�\��`�*�1;��j�Wm�����U(6@e�U�0��ZOmfDf��fgg������#�z/��c�V�].��	�҄	��h��lS]؄�b,�����9y�*����3�/%Ezf�h& 4�|���+�<�v��_K��� .'��v(�2�"2���eR@Ũ Ce��14�͢[���;]9գ0;'xho������:��������x(�4fUn���j����-Sggg(9T:Iի
�QeLmm-5��\p�����d�� M{���	b>��]�9��<Pu �T��ǥ�c��@Ȟ��A l��$��1Pq�M`|�I�����L�R�����к���F�U��Gt
*��:��Uĭ=�hk[J)+:�W���Ⴌ��v���#��f:���a�m��ƒ��.W��~�h8��j��%��y�J��[�P�\(k�p���]����K�h}�fC��2&e��QK��m
��A>Z��k^�`�M����C�'��Z�^�>BM[ۼ2����4�4q��О҂CyMM�������[�/3ݾ-Dx��'�a<P>r(��?~\s�P	(��B�CCCT˝�v���κi�$��F1ݙl�?��秪����"ch``$^�ZB`��
j��� #77`�Νn�4����~�?_��v����̵��� �==N�>��ֆ���&~Qߠ��`����+n�����"�W�� ���r��5*�eZkL�C��!�â0y��.�d|���h��R��Y�_������� �Q�V��J�qE�������Y�*��"��s�C'���~��U�H�C��*�W� n]eu�ǥ���hXI/(P� �}|n��dK_�r���u�sۋ�8��]�z��NE`#ж��L��j��������2���<=!65|��y��wd��PH�8<Tx	�څ�{���'x�6����}��!�×P^�tT�w��M��Ha�%+�פT?��搛i��6��7��_�1`0�j��x�����6_jλ�>?�#��k�(�/3��]��{���FO�Ӫ>Y��<��vc}G6l�G��0�J-#s���X��w��?�}�\C��iK��\L�Er���i�%e�>ǐ�2ұo0��_�S�̞t`��gA�J��H%n�E�TЁS�N4T�*��a�@�k Q�o��N��11��Y��񖆖�k�����AfS��iN󤜙!�xU��_�a^fІBf{(�x���F��5�����X�ɦ���x�u�E�69�&�KF�[���y�9]JS�u���1~r��1Ẇ,�v�I_n�jg�O?2~-��;�5���}����U�>i
�6�պb���D�;�z�UA�˹�sf��I���?&Z,�6����y�b�3?��[�~ H>yu�;�MI����y�(�}��Q�k����)�NI@���4�,��г�������<��s�I��p�x��ICp���>��������A��ar��c��C"�0FgA�ѕ�D=�*�/��H��>R-XL^;?���8�[q�'��R��~N��~$j��9�_6o��<�"���a+5V.���-?IB��_Ŵ��"z�=������t<��Ϙ����N]��(��V ok�/ū�"B�&����Z?�m��g�jJ ?��ǽ'@q�<��Hc�3��m+���y��fL�C[��rx�T�yʚ%z#Sz��3����1�^fp�o�=p(\xӐ@��G�Y�$n�!��`��9CF�u���~]* $mHtt�y�5���e���h1�f�\��l�8�v��ȹ����S��Y�p�}��KT��I��qDk��D�m4?bjا�<_��������ע�Q_G4Z��Q���s�[I��S|m嚆�>��w���Nk�J�[kf�]��D��PѸV߯��IL��P��D���QjҜ��z.�Vh��UuY�'��TB�hR;�ghC��E�젇dǻO W�Oga�z��F��lV(��c4DZnqM�:��oXD�~�ǒ��+��Ъ����y��*�W���GU��mu!Ӣ��]1�/���|�f��b���w�Y:qx7�+�NR����{
���LU�QZPO���f7���^	�y<[+O�b����zy7�z�|1�U6�bE'�G֜_V�/>r�����m��y�y���qc����L7�� ���j1T?���]�{�ȯޢ�1J�1W�� v�a^u2�^�Z�%}��k̖i:_��}ON<|���B�Z������8��z���c�:GQ�]�e�Nt���O:�
�Zk5�T���_�{�u����[��\�IةG?�b�4�	��δ082X��Թq�zn� �t�����^�ӂ]ب����=<��꣮��sng�|�(�D�'�Tb� QT�ۿ����\E}�U��S���,�� ������3=L$XP�<����'_����RĨ�t�Ǯ��*>��T���|]�[@��Bh���c_A>D}��]	�ˡ;�:D|a�(r��������|�G�A�h ������\*Z6�ˊfLJ�1�I$Uл�����+#]Ӡ��EK���'j$Ga0�7�Ȝ���+ оta8��l�fP��%�$�˃�ٳ�����zk��?gV��Q�zN��R�|x{�GS�)]J����@����[QI_���z�?���e�H�>7���!��k��(0�Bz�'��?-���/?,>[ܣP�>5�~楿��J }��-!,~�oϓ���NI�r��O}Y���aS���Yk�?m���O]0���g�����Z�&>`\�e4��C����W��~��<�w@���T��z�$y�G�⨵p�̀gj<��ǻ�B�l�Wg��5��&b03��jk��i���#��	>VS�'� �go����&vb�m�Wy� �C������WF���ܯ�h���QN�7����2�%�l���hМ&Q�,R�b���z��v�OL�G�vJE{O9�2&ND��j�"r3����~>��H���^{7�j���^���Pw����:HBП ����������8�`t�vA���/�Gw�B80#\�B�^p�3;u�[�ߨ͠#0�~H���z�Y�B��*l��h���$��Z'vdr�9NA��#�z��\q�$����a�p-��u�G:$���F�)���[�,�0��h�ӄ����ux%�+���w�k�A�OSXh`;�eq|��/���c#q�������W�g�d�S;���3��i8�.��n��jY�}b�)B�b��Ӿ�U����ζ�"��4�7�_�eIO+���E|
<d����לG�EO��5�#�����ݖ�^p�}e@��Qc�
>�;q������ω�tI����D��xi|�Wʀ`D�ԎA:���?F�fi�|d�}O�&4}�<u5�ͯ���� �S@m�R�Z������K�_~ =�(���4�J&x�1�Cs���"O�n޼s��HPr���1��p:��t��6/8k��b��/9~�l:�D���k؋;��7FPK�#��wB�T�p�3�nn����`��%�e�sLa'�8�Ϝ�`�+��b�r���4�A�If������[���,B������ݡh�է*£���ܦ��ϖӕ�����>;�u&=��ԙ����D%���M�v���o���G������_8҅��y&�}����-/���؇�O��MZ�F?�dk-;c
�_��.S{�|���=?�
5�Dǫ���u|v����v��(ce���p���0�/��a?JL�����J�6e,�<f��Ӛ�nT�O�x�{5�6~.-����o��d���B����4=(w7ۍb�-
�*E?�Y��|O0���V�+t���*1!��]�O
]�ʈދ�)��aޙ�V�]Jo��z�����75_���l��}�3�N�D"�Wv>_��0&�B�P6�g�����<90$�%�2D�R
�5!/p�H^
�3����|�S�����3����LMer�	�q�k�_�]Q~�2۩1�����k�9�g00��eb�g��l+ѧX��_�MBmt�AT�힏G�.�K����?V�n9>:3s���^cV.�禾8�w���>:zo��#�i�����0�3����_��H���U�t�9�����['>G�\���Ύ����K�{鳋x��.[�GnܦV��ic7�Q����3h�+oB�H��t |�m	>%j<�v�k�ve���x�[�������|ܲ�n}��-��5#U�~�K5C!��9�ش9����;�y�=z����L�u좍SAQ�--�EA�Q���0�J�?n�u��9��Ao`t4=�3%�q�8�%j�@�x$�*�g]i-ͭxZ��������pƩ����������"�݌���&5Ra�dN�[B����Fu�I�o��]R���VfX,̸z�Oji��oڭ�h�-r��|��"�s�����}�E����B��~4��3EcϽ�s_��\���{
ҚB�W�D����ϴ
�/
y2x�IΧG�K��j�3��Jta�Q�^M3�6�u���q�("��P�n�����-M5�%�6�˷�&?韙�ĽҞ�|�;��ׯ�5T����2�u�P��ݷ��Ԯ=�t[����X��V��_o�� _.ճI_w�^��Y=M�PU�e��������QHu�Px�>BQ-t0�"�����9rYZw�4��oThWI��ʼO�Bg~9O�77��n8暵~>_��L���nf}��SQ���^UXK�z��κ������{�dɦ�;Qj�	��m�F�C{U�~J�/m������IEtl���3����6�k�/7(�����Q-q�i���TZW+e��"Km|�]�΅�窅[�߭�c�x����=ףlvn�Ĝ��+=rc]�Lea���6F�g"'���/���
U�o�V���ی�g��z8�RN�v�`*�A.�,��j[L^�͔Xg_''L��xmv�i;Ayb�α��CѦ���q�[
&�żQ���8n�pt/��[��o���I�؁������w�����/���Q���1e�]=z��D��:�#������5��j���~\W<j#"���4!�_$�����[B?�{�c����'�y�V�<h�µ?Ͻ�����Ҽ�	���G�<�;r�q��7��������y/�<�>+�wm�R�-��F{<��u���$ò�e(���Vvu��� �v>�z��Οq��� �}빷�	$��DsR]�5�kb�y ���w��$w���,\]�d���ov�e;a7I%n�,�����2�Eƴ��x���	J.Ҏ 7�Rv&e�	��V�����G�S�ۺ�j�� !��,�xg�?�� �<1�����FFTM���褍�h���?|�����a��.�%�ݕ�F�M�\�R�c��h�����}1v��͌v%{��9n�E�!�͑���F1O�b=�_�E���˻݂^mb���߭psY-�%�pVAF�n�}վ?t���кGuv����9n�gr��e���<�Ke�M�g�(�<o�uվ�e�d1�FU�F�w�+���#k��#�cx�c�O�vo�ޯg����w �R�FD+~��/��{�	4�Kr��:�=��8�Y�s�gB��5�3��EO�Uj�},o^:c�{����N�$���k~&����xDA�'�Fn����M��S#�����Ky�#��V?N�+�B[Ԏ����"rt�`ZB׶�Ү<H4*�!���.�p�i��V.��l����T��g:48�~�2d�K��%o8�2���;qDe�ly��3������g�6�����JK�2w;7�D2P��Z��c����v��w�����D#���8�`=y@7�66�8��5$HN��!rA������]�`�`�%���73| �*n���@Ӭˤ��Ye��.7��?����h�1�����`�>�h��ے�Ͻ��K>K�<#�=N�C���O�a�J��[&f��(��,�ן*���2ɚp%I��1n�P{��6�U7;��R��.�}���d�?��7~�x�#P8�q�м`goY��~g��y�(��.���:�k�d�%���:X� �7�t�ZO&�)�'��/׽8r�8��t���6G�7�`���Xx�}NQ�,;X��!���lg���8�������٣����������S��4[��Qr��nK}��_3ދ��t�P���y���RΣ�#hr"8���]�������wul�>�4�f��.y�X��} ��{XRY��+�\�g�RY�Ԗ�a���Vr���	0<_W�]�ʒO��`ҩp��{�l��z�����llP��SR
���$�S?��W�w�����_��k�f���������Y��FܳepZ��AK�B}�5��t�YCN��%+�ym0�wq�m�*rnntWXXNrV�r�y���gI.nK)�U���d�,��
+m�z��=�GYH.	w��,X�S��$H3}�i݊�l���a
������Yƀ� {_�j�I���&��X�Y��x�����C��t�
)e�sc������խ��O�i<���	2���B��}��;7{�Q�6����v��څ��X��p�O��eGK�8R�<@��ѕXҙ�x�\�5���F��M}z�hƊ��-Yy�;=��TT<b���ե����j+��w\Qb� ̪� �=�7�w��6O}��G�]�3��}`a��$��`���,.tz������jֹ9߃zʼ6�ny��-���(ZSÅ��|��t��Ҧ#]����u{��l��5R#��7�3�7_���֭G<������Q9�n�-�V�b��)6�(҆��E|�|�^����붠rO���D櫻��7T*di:��M����,�����ſ��z�
(�x�AcK櫢�	��屟n~S>�j�7����cO�s㴶 ����Hi���v4O�;����[Y��`�f�-���6v��mvqjЇ�]��N�P�
� Ɵъҡ.�ع�d�dS8�'�g�#n��ir���h"�c�Y訲z�O�崁�ŀ���x�B]�������8\Y�"�:n[aa�mr�·���2~M��z(��ad�-���Ɠ��K��>2���������@Muk�Q���"M@DD���H��.�D���+��ދT� �t��Ѓ 5t����+��L�q���Ե����Dq���w�����f�͗���ML�L���� �b6_�}r)��ܼ�$i���Z�`{�&�>�2���V6��a*1mX�������-��V����}}9Rk�c ���~�M&���>@D`^�����S% _�����۾D�@g˿���6��`��o�^nn��m�<,Z��֧�fl�Qyfl���_+ALfj�6AɾP��-@� %�Vv�r�jv�]�0����Oh;~2�w�K�������uT�Y��6��}��qz�3X"
̼�_��+������<��k)�.׍�[߉��31�49[x-�����z@��%Ǜ3O,����>���c����n̾�)�e9R����l���1�"��u��ý ����,}����8������~��~dyv�ϢH���0�i@z/.0\��`/�t��WK�/�ڃFSd]� ��=?/��j��)'�J"������|4�1G N�1�8sȎd�������0����֤Sf[������,�bF>P�Q�m�t���E�_���1M��"@N权7�S��SR��Wm�ͭ����¯E�*����6;!a�w �����RF�Vğ]Za�
�&Eb]�Xaez��P��h����b�f���Y�����\y!���RU����R���D��n��d�OI�4��ծ�5ԍL���O7��8��nVy�=TI.�������O������)$����>	bylK�`}b�ȶ1k�#Y����	�>�Gg�n)���
���[?B�d��9������DgZ���D��?X(3�j����8��D��r���ݯ���LrpxU����!q��	b7�?��]jϠ]��V����E��G�~����˲D��JA��O����8��4GJx�_��V1F���[f��A���k[F� 	�G_4�S�--�.���+O����ٴ�S~g�%�Cς����@�����Y�����M�1�%F3���M<��W+DP%Z�����m���G"
&Dg��E��"���<��/˄sI�w�<�Iv!�?8���Oc�r5p$P9�겙�u(Тq�P��\N_���cd_p��:��:ъ�ݳ��;�r����8�s�Z�����R0�۝(W�������%k#������x�Ji}������Yb�x�+����3门5���o�j5���{�F�ub���A��V(����g���T��yfq����tt��^�A��#l����~�����z���Ϭ9	�n��
�"t���Qx�{ߣ����l��m��H=�w�#9z�����C�wD�)�|����ʼ�;��_�����1���Y��I�m�9$��|뾓׮olp����f��X �@r6�nI>w��¥*9o2�|����SN���jE���n�c-t�gX� ��F�l�1�o�i��6�u��6�m*�.��� ��"���ٹm������g���෈�<�k�ȝ7��P���Nz^�2�0(Ϙ�z�/�����ḅ�#pbӺ����/Ï�h$��>Nu�O��*���d��K�$�uüp��S�3;gm�-5S%��{;��G��䊱q�,%ƺQ,l�^��ϙ��\�f�~����e�q&����j{������zM](*�!AD��k�@e]����]�Ѿ�׶��?�ߘp�9#[�C�]��.-iSd��}�T�s���9���o�fFeD��Z�V	������oǕQڙ=����q�o�����<�	1ŐI�d/�VP��jS�Wո�r�F%l��z��/�%,�w�c�Ր�N��ON�pO���>���t5I�ɵ� 6�W�J`��6��]I���3�5�����-�צ�XA����2���?H§�����?r�]���j�@皘/��F��9]�]/�)c��'E�e޳,�\��`! ��J��x���ڸO���N_]��W=�8�S�.
�BT�\����<�������W�d�^~녺ףGWՔ1�w!n��$�aP��'yT���;$l��)g+mF����;sy�Dl���r�o*���uA�;ux��(�w���A�����"@a���	0ϭ������ ��e������g4�L� sTR�A|�	P�V�J[bzL����{�5+LzF�~�]�!�<N�I4T�'��l_v��	�;w�����%J}͌O�tܦ��w �� ?��+9gEe�@�A#wq���3�%
 zG�0C:���L�ē�|��+'Zl�KEتMV'��B����1Q�?P̯=�^�R<��V�>	��	��\��ܿ��8���"�vy���� ��Xw�#FT�J�?Ȅk߁55�J���r6h��Ђ��<��_�L_M��Q7Q���]�4��I]����6G
��!�%�N�0�ĩ�|��.����3��E�e
�`�R��31?��P0� �mAP�t��	+oA���I�mQJ&�����^uf�Y<����C�.. ,GW,Ӷ���-a���?��n�Q��]�buS��c��\�N]���1��0-����}�-gD]��4^��=�BV�uR�C��u��'؜\��z��YC�F~�K
0�d���X�6�67-��D9v�`8�<�k�KF�Z�{�7H1��k��ű�#�Ό=.�.!�$L�����'�:����ME�Q����ɲ�낕"���/��FD���.�(�1�V/1PFU�ץ��z��'�2(�`��MY㎝WG�OO�ț�1%��V�*�
��;V������fA�TP�$ى6ޙf ��`5ۄ��(��k�җ�9:� �/M���:=?J���ʵ!���B.�S��b/��f8� S؏Dw�pIW���?���7�sf"ց�`��`�\~����?c�ھ�Z�� ��P�r[Ɠ0G��M/�|��.�LY����=r��~���B�jN��*��A1RDN���*!h��&�`U�w�Km��& �&����1�D�+�V��/�X��NLg�r��֮�����Փ�͘���.
#����w`(� !�#��h)!�u>��&%�CZ'�<�Zk �Kr���It���C��h���N����eމl�&¡7�)V�n2�\D x7�41�`� �
MӀ����T��q�m��Aݐ��g`P��l�˺���}u�������U��'je�/L�]�p#I��͛el�=��hB4eY��[Vji��7�(S�%Ǻ�y!��U��,&�ƚ��|��@����[�������	���E�G��!Y�唇@��|T�>@k�L�z}3����aT�F���$��!�DP3���<q�^���.�oߕ�١��%w2�����z]*��3^��jw͞��2����=��N���h}X� ^�T�_��Yk�<��V~�bt=B����G����.a�Q���a�nģ��IH�.K��w�Y���s����E;�MEO�x���M��e[�R�>wc7��� g��&�����$8&*h,��ZoՎn".���m>�v�����Ug0��VK�nd�A��B��onv����-��sL�y�����η�
$C���C)F��W6�֕^����㱪�x�`�@F�m1���c��V6Ѭ�6||�}ϱ�K[Q�Ǿ�7����G�A{'��ktCf��{��� %���גվ��6�/H«P�3�����f�������79�@D��A̯*�_����ei`~c+���9���}�_2��u���˯~�IdÀj��טq���Z7����r=�[O���@Vht�u����&�8,���ϻ����C�m��Q_����0�3e��ru���+�~��P	y���E�i����l?�.�+e��g�Pa��v��j����2�Z�>`ҽa�hFJ�U�=��vР��K`�1I�48���8��v[ru�хL]�>�/��I�c9Z�`>r�j� �re������!��~��Є�09@��uC�a h��r�3�MgC�P0rE�r�H3t�ָEVT�vP���;fB�������Y����{|��z�u溪MHK費q�d�p.i������ʥ`��q1?b�*<��Z��o�����z��M��A�2uaJ�O�;�==�*�'��Ӭ��5��aKKߥ�ї����S�c�5.�����Փ��a��F���Ȭ΀R�����<ն��
�1BXHCH!
�9_�s ���sJJ}�O���JD��]���h2�9<s�J x����#2*�YD�2r�W塡t�VS�bba��DN�tsJ���ص���R�Ŀ���C�2�r�P`�I����AeE3��`�M��S��ԧ*�����z�D ��MJ�|�E<I"�i0A++r�I>nb�W`��;tA�L��u|���]��͡�⤝aȟv>�Ēg���S~��v�&�'���}r�n鏌�R����-��\�xRmh�����)��_����56G�L�-�7vح��C:���Lr`��K�J��5����OV��v���C�δ�f�3ej�������}b��3A����`ѩwŐ���R���T�S�6��MzԪ��Bb�va���%_�h����8B����ʤ�%v��)jhZ�������bb�zU<����P��0�]֎i��ee��+�y�c�un(ĸop�6�����:|�fw�'M�@}Vhܡ�Ս��a5�vW����M�%�{�=�%�������k��c�����|�W�p�����<U�����!ccf@�=i�Ӓ-!�;�?)z���[��V�?�G^����3���^�e�U��ۀ�B�0���U4j��j��^�0�5E�_�z���G�{����Ժ#K�tj� ���֑�.��c*qP���9��È���=+�:9�D �ȴ9_�ȴ�j(�����nMvhY�FN�V�6�/��sy��~3O_-�_�ڛqΘ]Z
AL�pwv��s���+�`�C �r��G�^��׍	�l��('կ�\6s��F�vj'��,�4�jT0��$\���b'�묖ҷ��?���m@/z}I�Fi4E�,G��V�.0$��C����ϛ0u�����6r�n�6Os��/U��"~x�ă��������Vp���MI���,\��Y&��:�&��C=�K����^ӧ�����@��+�4q�&����t����\ \��+Z�У�w��*�.��g����>�5m�N��k!b�o��:aM��lc��$@*����y��C��3��$���㜍���Vٞ��m���W�z�p���K�LV��s�{��'�&V�=� 6J���Jh��g(��/Y�"���	���N.��%Ѹ�
���m�`J��-\�<�`t�i���m�'�����'/�Yg���MȾʆ�פ�l�����Ax����b�X$|ʩ����d~0�Q��H]��j�i� af�"��ѹ�n�h���ݬ�M�A�w�&�C6.�4].ГX�5�ĥ�z�$�S�)��6�0�+A��O�Ϊz�c�j¥�Ϧ)�z�3���
�4�`t�r��7���SH��0����zD��V�2�����=��˥���]�R`ͱ�O���[�%�-5�E�{}%�Rð0����V`uB�z_nO��\��۷�Ć��>�"7[��;ۯ�K�{@\s���}w��7��w�y�k��O��/+b�s�W6���':����cx'z�)>�}�jpֳ-�%�Y^�`0�Q��<�@ �iZF��'sD��O�������L�B{���\��Ç�ԓ���~��7��SS����*���CK�w�]1�X�s��͕��L���Cױ�.\��LP���Þ���Ui���R�����M��ğS�ֵN�g�oکK��̘��ж��AڊW�{\����K��B���b��


�^U��?��wWޑN,�.�[`>.EY�Ӌ�$���'��C�S6M ���ͧ���#�@_�D���wS�$'m
[�F?q@W�39�Zr�뛝��o_��U��WL��V��^-O3���,-��ګﶗY^>Ї��;���,�u��%ꍤp�����z��yz�'�8�h����â��_k��ը$!�s�O���S7ט��966��f{�����/�x-�wq'������(nܣ#Z���M�E�5�GВ)QS����ᮙ�����h/y0p�Q�IȺz�t��b'���r_���Z��_X��3���}]�QÿӴF��c�;��ޱ'.�#�tu��P����̰�ML|,�b�c��5����p�{i�x����rH)R w�mz���q(�	�ső��������P������-�:=qZ=�[���T�>5�8�-�)y_�BA����8��`#���7�(<�x�V��4�|V7��؝<Y���M	D����Rt�ZZ���n��4xȠ�	���b�H��_f�E��k��L��.s�3�tl���?.�u���a�z�|H���$ 6m`/������u43_5t=
݋���4���O�r��&���`��s1ȰDጧ���~� ^�h�3�u����mΤ�g��y�4R��K�154-�уc���y�n�p���J��Ŏ� b(�{��l������9�#�}9���L��Zf#����D#R���`����p��r�Zf6~uh��7�/���&E���`��.@hy��}/��K��竂����ٴ��.��74�I��7N8�O<N��[|���>��'�y��W��[L�D��ۭ����l�]$� �9@HbD}�2|
��)S���Nܟ��<o�y��cʰ�X�~��W�l�w���n���+4;�k��܀�=d�V���,kA���-���N܏x@zl�6��B�˫��
�ߊK���������g��i�I=���зG�q��n���K���P�575��D]Y"�A+���,�)R�lj�����Z|�,M�N�|����]�魀���N�$ǌ0�7p#n,9�i�Ue�;t¨�3�ܐ*�Gp��q��HF��Wf�J�H�U׳��#�RmF~��4F3c�?B�iq#�[�p��hϔ�{%4�+<���C���Ӏ�婶� 63m��3���G���I.
o��q
$tu��^�ڳV4)�:9�J�M�z�\�d�f�I�˿�be�oi)2=Z�LqM�Z>$�d_/x�'��s#���	�� WKe�������p��feQB�� |��͛ae���&$@���q�>|��U�@~��h���pY��ѿx�A�č�n�]�4��Z��g2튶/3�'��m��y�����ڞ�H@�:W��H�8�-;X�͓jXc=�d�&	
�ΖO��[���Q��y�o�hm����Q �$̾P}g�Z�Gf21����'��G����J�4T@� �2@�_8���n'5��:��g8@9�T�-}]Q6�a�ú���9��!`���"�W%!����4%��8PrßR�r�p�(�&�T���')�+ޙ�u���Ra��7���D/1vm~��C�pF?�h�Ko�V"m����FI�QBC{_��f�B@p+�(��縗f� {��T^�[�7�R]�Ӻ�|!9P�:t���l<썥��"��'���@$K%��E�6�Ѵ_�L,��Z��b8ߏJ͏,�H��bx����������z��O�u��!��MoFC�A�<�*��-���-Q���!�!؄�^�$88����e�F�^������3;��2��"�j�#�h��n! -�6�����Ҙ<�T�&���U�_R��F�Q���I�n�7��Y: ������O�7@z���IP9�B���)�d���v�g��#�ݢ�2����3��g��a�?$KQ���+E&��Hv-��H6���2v�Z\a�����ˍ��ɝU�c}Y����G��%��BuW7��a�����#�B�ӟw���F	�x����i��x�46�Ok�:1[b�\|?���_�)e�2vy�C���v�_��.��~B&��J:�^���o�k�0H�3��Df1\���O���&֢r���s�v5����M�D(E�?���:��o�+B�`G��e��Uw+��R �����v��'�{�Lq�*�qm;ZS2�z�v�G��ޱ|I��i�k��h�/��"_�3�/��.�Ś0�W���h�T���r|��Q���;���D�����{6Jw�-4���S����¡��a�@g�SIؙMx�	����4� �^��Ӧ?EFl���4����V����s8_�SƑ:���7	!hty��]� �z$s2�>{��i��iK݇����'
=����~` Ȁ��;VIL F���V�-��ȿ���P������ˇ��W*s���X���A�>��p�R&׼��,��x���On�d��XPl���͵=꠺�;tKշ�fꞀgh̠Vh-�WЉ'���A�R!*��$���" q#�Ku9��Sb�2�Kc�0�h'�D�j��MG���h�0�
�pI��M@֝k�z��0�3Ҙ��<O��x:�����F�}bk�2;�%����a[��B�=���]`��r}�H�9�׭:s��Au�
�+j��wY��$�-�ftZWȳ�l�l�z"���A\�{m
}��C�&|w�Pv�V+t{\� �v�{x'</��I�bh�'��ۮ�q�����ա�D��w�m��J�8���L� ��ee�R���h�ݽ�Q;�M�0哺T4|�N���c��+�U4�b�,"�ZYJg�n���V��H��Nz�,��$�cx�W��zl���u��*4�c�����v^��� d.9�D���QqOχH�N��N��+rQ���n�����C�����\p�(��G� a������۞�3+h�$�ޱD�?�9���.#�5�����۞fKV,�����o[�U;wI��.���03�4���EE}pYѦ��ވ�Ҡ=������y{�6F9����D��3`��ZK��s���Nh!���k�Mȯ\�#ψ~��̊�:<�* ��e�_�_�@2Q��*%��lΑoS,�4��(55��_�e���P�=R�ϓ�0V�/�A�G�0aM�V]�}���vv�_Ǆ��X]�!�a;|�P�v+f ��*Se#��0��W(�ԟoTi&{<J�����%��2�m����_,Z�{�)��Q]��H�qA����#�4���C�<����`����3�P9��Sf��-2l��U1t��2Oխ��ئ����>�	\���i�1l,�-�G2� z:���K�b�(�g/�ͽ]e�k�V�o����߇�X�5[D*Ĕ�r3l^���ajሗ.2�}��k������*����}�a��]����DG�>A~�i �=��G�l;�s��,݌�\��	��{�d���{�6a��߁g��f�����:���@��6S\2�"c�QU��\�K�Cz����� Z�q\/��}P�R�{#�{�N�}b��\�;pxMN%�Z]U�;�MՔ=Mǵ�T�~�W*���4R�h�@��4Tp��eWC|�Z����̧.	Ե>I
�ys��9(�\��>$S���[t��l�}N�t�lD��1�p�⾖{�i'#b��D!��w��u�ڑ�ܢz����J�Of]i���'�5��.�7��t�1)$$�/���9\b,�Ю�<��R�ͷ�x���32�Ӥ�ě̈s�����3��/P!���Pڽ,,`j�Y����E�Y����ס��r}���3{�C�mz{� �����FQq�&�Bv�Lޚ^�v&jz�;bί��f��s�9�j|���9��j��-�k8��+ڟ'F3����Z�;��O��@�Y�l�8I:�4�`�-}h����(���s����M5�֓�;��UJ�Y�h��_��=�Ϋ��&��z�rɐ�ce�u�I�YO�3��o�p�����&}�&L%ת�ҥm��cL�,nF�� ��rJ�шG�e?}r��@����NL�P�V��}ݓ��U�%z�?�09�e`�]� ���ȿ���t����('k�c=��K�����9^j���O�'�L��v>�}\ڌn����h�y��ٿ$|�gCo�WW���3&�J<}w���߄]1���U>�����TTCe���Qf��C_��^�5�в��L���e��XD���#��c+����$��З���=�����m>d��~"���\lzQ���`����SC��ܕ0��-)��G^ooW�SN�}|�����Aq$�.4��o�'�������T��vy]�p4[n�����.�us��D�E_�C�G�<X���iV��<��C�U.!�@ٰ�7sj�w���)wؽ92�mPr��v��#�p>.Ƞ�snæ<h<�_}�kʂ$W˿��2�!h~����IR>�}�2�$���drа����6xs��Kx�믁�;˟a����2=���%���.N(Z7�7K^��I��RV��A��8XF�����;�:�$9*�宷�x�iqtG����뮛�)��*)��{u�e�9!���!���45�ﾎo��H���bN$n����4�Y���q0�v���A�Z��ס��&J֤�[.��x���V�ߠ�gȮ=ݭ���m@���{H��,+8VX뒞������2I\=dZ�C�.-��giY�<x�W�T{���9�3�*Z��܎om�ѧh]��:�"��;��l�ə��\^��؏}{O!�p����*�y��VQđ�L�����s��t�m�̎s��1q�>GM�+y����F����_847�آN�HR�%���F����D%B�Kd;��2�����`خ���fbe�JY@�q�toL�|��	��j�����p�J�G����o�#d�u���Q���^3Z�@��Ϝ��U\��ncgș�!=p'�@��˂�=1�D� �qK�\���)�@g+͞���;�I�*p���X	?��#Q���f�m2(r��4�|�'�DT�y/����AIթ,��xX�f�`�0��� As�jd0p�H[�cPިe@����Ĥ.���5Ѐ�y
�X`�n�w��*��w8Q��v�^�F�M@���]��R��
���;;]i�E1]��K�n�ȇ���sX�^>oS��5+�]��ӝ�s�
�w4�x�6G��l6楦`�|�[	��V��s3��C�Wj��A��^�=ً���[P@6��Z�1si���ېk_��Am�����65M��6��	�J}ͺĊ���>_|�sL���o{�5��a��,N+�+�^�t��.dj��-���%�C���d�9����Q�F��?�,��/��-�+ۻ�{G{i�"F�J� =��"��і�<����0|A���r���7m��;\>5��l9
]z��&g��7?I��$����JK�s�����.�����it=��F��޽w��{�M.��� �̏;��$ͼ҂O0W�����pE-��2"m�����l \�ں��JW�3�l���هga�8�aE.~������XQ�#�V�Y�v��.,�6^�֕d��)�b�<u>H�,}۝�xf�TY��+��T{7�.��2Y�mw��oy� u>��tjyѫ������tM��#��&���wK0u5�d�D��<_��T2��l�}b���6��]�b���3wl�?��&���m����Q�Ha<��5zHrrv28亡�:|)�
$��:)2ć��t�ŅY	U��G$`�R��c��k�?S黆�RlW��g=��W��fӓ��dҾJ3�Ȝ��͇����L�ȓ��T󋈣��YR���Ǭ�K��F�C%dOS��a�e>QH�8.�|*�uN;*~hD��K��y�+����t�v�^��U{�l}{l���f%�MŅ�*{���c���U�ߊLn�Nz��)���y��#�1����:Ol�nI�Lm��3�G�"
,�i����=\�S�x{u��cJ�b('�q�Y��ug���V&6��1��y�!~�t�o��2����'��z4ݘa�+����\���	��J�vu�1��Nyɨ�xl�If�\�ע��KS�
D"�j;��c��}o�"��C˙�����/{�x���~f�'Mu����L�N�$X��iU"�k6q�in�����d��B�dt������PZp8qߐ�`�+�1R��L��RD��qj����&<����}������nh`eկ!��u�z�
daeW��	-�������(>{":*�ֺ�ʦx������,^	6���~ɴ�'}��	�����I�r�;��p%d#V����/<k�8�W�]Ȑɇ���Ϧe�Ad0%�f�Y ��D������c�*���w:�J�ߤ�*k��{Y-]X0H[�k������x��{�J-
��m�O5^,�:b�M�N�W�����Xi�Y��\����w�K�1� ���ɘ�~RǞ�г�C�\S#��uhE��7�d��F�γ-�b�zHD��[��&,��	�&k9|���N�:��n�cռ?�[�;�  �G��u G՚F>�V'�53�,^`9uR�-�\k@G]�3��Vvamhv�j�w?w�c�av!]B����0��ǚp��O0m������=�4���6���}�|����.�+�tl���z_<uР"�JL�/%���O�]������������xJʱ�����/�A!`�I~�c��0�� )��?��g:��AUV�)b���](���JtK��|xF�iu���|��i�+K�{�K��z�v>|9&(�y�Mw��F3�r椷S�6�fӃ^
=���]��AH�=�]�w��^������ٙ�#?�;��R�ΛWs�-��Z��X��.�e��4	Z���KX5ׁ\f�0�P�'��o�wp.�+��)��p�H�OqZ�ܞ^��o��S����7���})[)�� 띦�՜��u�:��.W�5�㢾���C���Xn?s	J�������d�fއN�Oz�́ۉƈ�6:α�V���c��t�8A|�&:;��^(�䛩8{-˱�X�x|i}�qs.���`~�t	/P�C�ޠ�*kll�&�K���IrY��_��V�*����,�gC*?;|;��$��\[9��g����%w�-3rf��RS�����\����nwWh `�����<jqјzg�;���Z<��3�Bu0�C�=9�.F�#�4����p���۸
�Szj�O���giD���AJ��z���q.;������
��:Vg��T,1�S���e<3c�97W����5�y_w��S¨F�G��c��bC�۱y|un�O�3�/gؘ!���8�A:E����崴�-9�p��-�C��"��;�ɧ�+r�b�O���&ú�E	,�o�	u �z�S�E �'~�n���u0g'���e��Dا�Q��w��a�)7��� rX~&�Ь�?�;�����4�x6���>�It��^�h8�z�RK�y��]�r �vF9�.�%}F1�IL�L���ћ|�_(��\E+v%� V�/���EF{�^AЮ�+wcm�|�~���5����3�V�sl���q�pcJ�).�b��Z�sK$�D�9=� ����U܊�N!K�D��?�������^B/ul+k�o�t�>����c�Y��͒fӗ����������k>�����˱��6�rR�ih�T<���+���T�o�Y;?�tF0XC:��xPC��R���gjs2��e�6�ɒۺ^o|��<��ڻ6ј��L:6����!��X�x~���5L�Ce��V*�m�'����1�nl��;�T"�����LZ�V�H��GQ��<�Ψ�����!��@#4&�r���y	������{'b'�f4rJkн@!�l�Iv  �+v�u�c������2.Jo���iD��k�9Bf�"�CR?rCՁ���n	;�E�Oy�үcz���w���!��z�։!��7�A3F�������y��K��x��l��;�ʐ���"��;��;��r�����~��Ր��f���d|���K[&�Уry�!����^���H�t��2K=I�=���G2wD�e��gg�e�;�G�-]���q��?1��X�����=��%��,9b^Y���9XE2kS?���#��������xI!����	�z��e=��TN�O�*��i@��)��U��c�a�����.&X��%6���æH�[7��V�dn.��U �8	�f	|=���Ϲ��ƪ��gGK���o5�ͫ�}����l�=�U�G�})���f3��k����p����OϾ��L)ra����묁�� ���� b*Ӿ��e�[M>�3�!�aGҤ�JH�#��چ��}�V�ڠ6���#M4��\xAXi�y�����V�*ȭ򘡬���� ʚz��XD��y����S��Vs�4�j��� h�~� w��Ք+c��b��2�����+�_eW,�ښ�g���B<k�^a��?;���3D�k*S���}.G>M��$D�����p�F$`~?;3 `��Y@�7\�[U��^���h�+<�����?��jR(ͦ�x�����	U�Ϙ�\���KM-$�^�o�Z	s	=7�bj/�;��>�k�͕�G�l*�U�r�#0�8�q1T8W���﫩3�xݞq�6��o~`��R%�t�3ᖄ�q�Q8�:����		�,�Z�L�&�����5��?�O��Á���=���WR,�p���be��tX���j g��K�\�U,�#,�f��s��Ba�%���vM�n��ڔTL�I��l*����!9�����P��и}-��8�~��
#��̺�#������sT��ʕM��%��8��NI7�D�����5"��v�coӘ4Xp��7Ph���5/�� �ć���2D(wW�2v[�KX��'�R�x|nm����7JF��)����s����|�y����>F�v��)���uc�klx���z!�Dl7��%-�Uͬe����v��yl��_��b�!TJ|T��.�E��M!b�S���rWO��+7�[�X�~&u�-n���q��6=�4h�<����Z�J��#2�'�	/m���B���oI�Ղ��G�b�����P�I6-�<L�}�*�)�f�@��ɝq`��ƀ��pb��i�աnV�7�f�,�$[��^��j�~@���^�0�#UYqB%X]M�����<ƨt!9�_q���'qrY$�����h���6��<Z�Z~!��e�!�� U���� ��Z��q_�5�{�Z�Hp�3�Y򀩒E�٨o�VGP���8P���[�J[>Mό�hy>i!tcsq��e û�o�iI���IG�n��R����C�U�p��&�*��襤�5^1v*���~vVy@$���/�4
9cT�uP��E��`�Zn%wQZ�B�X�N���ݘn�yX�|�������!�G�~�Ϥ�J�v����ٖ���ia�����E�%<�s�����~��3O�ҙ�v�V;����@�c���+�*�;M�nQV�	W ��5</�C�{�+��sI��V�s������C�S��j�>����T�w�v��f�L[OM���l�lt�*7˧��|���B=�p��}K�{�@�\Q��3��K^vr��|�p�[B".�����*��iU�شp,����%}�&g�N�9�U$����ݿ��z�+*(ڽ?L	G�<� 8��k�6��Su��I'���v��nO��{��YTԚ~D8��~�v�J��˾�������<��[S��iP �r�Q(����I�n!�:1C����V3�`ھ���R���F$����BMണ-����ĩ�;7#�χ�W]�JfM;���يf9��K��/a5�@��6��0	dLE�)M�O���囘Ҡ;�%���d�L�}ir5@�*ܦ^|�78wV���>�>�T����}���g=8Y?���B� �h����v>؆��9���
t���������V�3a![��1f������X�6..�A��J?��D�D�fP�Lw�价������{�u��%���dX�	�[�����Ý)�د-��e�{�ꄄ��b3I(�c7����+��n������a��-O��V���З���+���a���"	�L�@Oo��m!�]�o�^��n�V������E�rZ�UN�F��#N������ύ���CRa���)#]�����˙���=b�����۱��T��Mk���{萺:6�"B=�\��z��@�-1)I��%��|�����z��k��ge��q��qҵ�Gb�{KwW�y���6�qxz�I�I_���k:�tv��N�8U ��N�QլJ>y�z������e���pm|3�ZM��0�S���G�%8�����~a��G�Kv��):TS4<�	p�v�t�1�,�_�-���||�Oq�h{�ϛ�oԯm/�1K5�C6��)��!�Xh@�nT�?�=��_>��i�br��V �_��Yu�A�F�lOSs~��J]�|�ⓁdIm���"[ev�ߞm9�<��gO�S2U��5���KG�7 +	1%�R(���B]��~�-��S�<��G����t
�+$
��b�c\����ռR���AK�̈́n*�󮱵K�H|�Q�Y�s졹�.?�n� �R9��*�Oe9�N_��oB��?����B�Gf��x�'��w�~e$.��Ưlb��7��	^B��
J!�g��.L\xA�2ojatA��%��ʌ�\����i�I��������a`L�yNVtȘj�h��74Lc�O\ nA h�K��x�J��Ç� �D9��V�l'���Q�:�z{�U&�?3:q��W�?,0fA���M�����2�WQ@ֵmtgL6�`Cᮔ�(��� N�H��:�e�4T4�>n����>��F����[�P�A"��N���|�'���2�����wH���ϟ;1����Ӯ�ۛ���Y�g3y������I�� � Q=�[�gHstk��\93V�^s��T$���n�ɘ����
����%($T�#�(FW��F��r����T�-a8]Rs�ӻR:l{kވT�U�l�I�8k�M~ʞ* �~�dn�]��m�O�w�h����gtV��
l�ig]ñ&|��IK,���dM� ��}F����@�UP*ؔ������Sjj���rN���N�d�T��pW�O����*�5��c�â����QDP@JAR	�F��Α����D���ib�!��$��;��<�������>g����^{o�K�/ ��p�n�&#��;�V]w�����n�T�n��S��7�M�J�H5������նGo.1Z���?�C����~9_�:�TM-�d�H��$�m}�[J��
�z�Id�L��h��ni\s��d露 �m�.&��8Q�>��7����h�ꃜmY���C�����ӏ{xU��)Ȳ�I{E�󉽺��L�� QL�XwWn���F-�\�o�4K����2c��Z�5�i�,�T�kڳXJ1��F�C�[�&��C����֛��+�
�	��y}%�<t����k�R\\�^&b�0�v9�p��^� _��̒��KXf�[��a�.w�5k܎%O+y//�l�;�m�޵�"�U���W�FtJ)\��3��I��R �,	f���i��mޏ5��z)���t�Ҿ�����"&l�z�:5�\�(*�`�W�F����T?�SQx��Ӿyg@T��t�<.�l�dw�6I�+��:J'�۫�S�V�#����t����Ώ\�݁�o���&m�h����ó큣o��ioI^8"ޠ�q���#erfhRV�[K7u�v�H	�&��7a��j���lMJ~������y��̾�o=%A��q�]�^%�*�> �65=wy����SX|�f��=M/Î�-՜�@Hǟ�S�����ѣh���+�~&�g��~a����L�l'�����Z�L;�I�M54w���f���W�u<�Ϧ�t���pG�DW��o\x?�B�bO|��^J$����t}��4D���d�~�[�D�O����M�+��ۺr U��T���B-3���؎퇣g����۸�j����,`~��*�a�C�W����}���M�C �e��E��Tu��q~���W��v�A�I/̫P4���x���u�[o��K'��d�mC�����[X�NKb��V�_]�r��F��Q���1��cY�����Z4��8�/'��8�0����-Ѫ=DgMX��s������Pw��)@��"�Ï�؆�O��Ɔ*U958'[��o1�7*s�rbп�/��ر����Ľ#⟬8ԍ"ӝ:�_�����h$�u���ER������Z��^:'��}Ӟ��~�������[�7MI������y��n�����e��;r��F[����D+9ܓZ�FW+�b���^V�ֱ���|�8���>�z�k.�:΢�b��2�0i�;���H.�'�
-'v�N�j��Ή!�W��dw�����1�w|��-�����D%r�o���dp��_�'9�'�����"�M',8~iZ�,N�FQ-��w ��h�� �0X+�
ƥc���)�^$��N��l2���߸�������Jg�H-�9��#��i���~_�F����f������e	Q��v�ʭ�mh�r�5�3���EC���{�a�gktk��=�-�����L݂�`	�[5m���t�'e1�����l�F�*b������dJ���a�=-��M�Z}��2r輰��|�nw�Y�py���&>}��x�m��%����Al�B��z�O���t�L�B����i�nOm�Ƴx)��o@<BZ�3l�g�K�����W�򎄋O���G���� Q��5�਱C^����X?@���΅&�	�j�-"��C�m���t�FI�
�ĪK�͵�$ej������F����)��<U&��^�%SL�$��\�=���^֠�D�-�]�Xţ"-m���3��S�bه���G�8Ḽ�S�r����lި?;:b��7�.ǔz���3ti۔��?��=P7�}&n"�{fjPk�ݢ�\�E�v-i{�r�G�I��	���W��-�c�Ddp���^{�R�&]u���ˎ�K�!#<��Hɑ�-Ȓ�Ї�WuI�5��~z�f)ξ���� ȵ��n��I�/�/�K%'�ҕ%R�O-���a�+o���ŋ�h�ܱ��o~!���R�r(����h�y�S�{��b�P��+	f��Dv o��c��OW�qv�Ep\��[g�j���+�EF>���}��*��n�5�ۧwg���rw�>C:�VG�w']�F�ւ8Լ���� ��y張%���cn�2��F���@NA[�w"N5f҄_ԶT��,Mz{G2�-[���9�m^_l7z�{��.Q����g�+��̭��y�nL��Vх3��֧�9@���d0Mi�w��3��$گ�LH�d+Kˁ4L�g_J�}�4�˭pM�
����e緧�dBX\hr���u��"� ��Px�[j����6�R�7K@�2z��ܐ�l���Aa߳WEפyM��||����s��y��,�`.���H`�a;���&?R͸tOa�!,���6,�6�8�L�{�;�K�����o����U��c��$SY��}O���˩`�AR�{�������q15��W�H�J�Y�)j8Ơif	�ʅ�	�b>x�Y�P}T��֠CrG�Ϛu��~����qLx�,���
��}����v�j`�`Ũ[��G��qQ�ب`z��uӄ8����{e�@�K��]�.���M�����mvw�T8��SDJ=�I���xϷ�o�;����}�.4�|d�R�|�#L�:ܞ�(r�[�� �V$���g[���� �d�̽�W��d7@���4N~�|��&Цg6�A2PC6��� �q=#���E��� ����8��7��,Iz�>����q��X�t����/�T�1����I��Zf1�s�/�~����d�:���4���a�h�Sy�����Iyw�Mx}�U)Mf��Y�ԥ�?쭣�N�˕N#��v�/<Zo
����LoDtQ�p���X�QC|���ŷ�H�rJM~��#�;ـ}H�fJ��M�6����:&7þ���&���!(�n���������U��CR����h�O(-�r`���o��c�V�����D�өF��%�D�ʈl���n�s
cA	��6��8��:8�F�ܯ0�߱�q��!!�'-�wah�c��J��j��VV5�D᳐s���K��#A���=E��7��̻�7���-�$-��<;��w">�t�s'�	�q9����|��ӭ!�-���\c�']U��eG�pPs��\72�����N�P��I�v�����m$��k�|�_��G�T���TD*��*ؽ�0��T�JY_Zx�����:���j�L7��(�scaQ��k9Osvq!'����;<����.�m��fa
K�����)���C1B-���	ub|�p)X�hC��9Ŀ�r�8��`�j/g�����ظ\���s�Ol4������E����
��=��2��E8�Y:�cU8�&(�LK<�9���n7n�uç��X6�� �/�z����I=�`D�?/�]R�AOH+�օ!JyCe~�@���U�/0�Jd8p�Kg<<���Ϗݷ��ĽV"�>��J����&�L��Aiâ�gK���Oy{-I�	�w**��%i8��r_��Ⱦ8���K������tk)JGz�%:��۬C^�2��(h�U��kLh,��eY���ي0� �~��8\�dW�/Z��%���^s���~=,��(G����VUJ#{.�n�#;HZ���,�mt�	Δ�}q�I����3�@@�������}���Z�E wk^���2�H{��]W�6��iy�O�9��p���oZ)��-��ǵfP?�<n�տ]�$s#�Ȯ��q0�(�u�'�|����щz	x�j�)��x�x��S�?vj ������{d�Q��Sd�c6��x@_��Mg�	E�TZ%�~EeO��/d ���s�l@6fLa��������P̹G`�5����+l�B��0�/�B�߫1�VC\�ȸJe5|���)��faҲ�9a�S��\�*��F�JUW�e����9N�����$x�ӌ���%U��c��
��0�Y�����y&#���X�=['Bt��H'�-jf��4zI���f[�W[)���������U~�Y5�Fn�����#w)��C�B�Q���A3�h�|?8�%������ݽaӐ�K�?t�&Z��G�&�4W<����g�}a���@u� B�]EcjLC�C����H�D�R�+n��{�\���:E��9�m嬥&��!�Z��<�[u�{����$��}�Z�
�P��a�K�%��Z^�*��\V��/,`������z{ �����=����n�j����=�)�%�M��Vur�z1Kәrq��Y�OxĵR�!|7�'�� ց7�".~��T���-�$�;{�ȣ:d�`5z��h��MP��_�g��"$�U�X�S/�n�=^��j��j%�/��o�c�v�뼸4Nƒ)+=�E�A=��ba��|H��BM�Z�e�53d��S>�\ż���S�^�9Sw���#7��=%�F�<Q<aoۗ0�[2d@�M�$$4v"ė���k��R P�tϟ��ꁸ$_Z7��i���^h�k�nX�����I�I]������Ȼ��ֈ�ɰ_�;Y6��n�ʻ3����	\n����������1�\�e�Jq~���jB+�D���"{��
W���J��s��/������W�qBGme�Q��7W���u�Dp������p�Zf�P�N@y��3GY��A.q��T��q�%�����BM�]��j��ϫ�,�Y�F9�~v�y��l:4�M�t�b��_�=�(%������}`�������(�����T��q��2����G/��1��Wn��L'���jz�_�b�(9��3���/hH��q+�;Qx$J��O�&,\���Q��Ҩa��>����v��̢ח�s�:D��}D�x����.B%����l�Q}C{ ��d��C9����7A���K��8�)�z|
��)��d6�ۈ4�s��r���Y��ဓ�23����
9�3� b/��ǅ�1���l(��A�7�����L�F����k��z;��/Gg�x̣��?cbW��r���,zEkz��I��px/��]�5�$zM�F%� ����s�A���2���ez}ݜX{m��K(\���?�0�'�}�f.29��.\8��U�\=c4ut�T�c�0j��x����X��U��
��=�AT�@���c���[��"ݬ��M�0T�4b���]I^�K�nS�?�0���cN���a4V\ӏkT��UŖ�oЂ��㷍����,�����S��=ψ�r�N/#9'����3Z����d5�I��
���W���[?��PXC{�:r,a�R����"�Na3yQum�{�b�\�)�B�x9�z,=7�T7�KNp�JDbb��b�x�洰�����vD�#���B�V�8�6�À��[a� I�kq����;k�gQ���ۏىhO���;��:��ɨĿ�S+��`àQ@*�ߚ�EtǗF���n����{L�AD���[a��"�o	O[�/ �o�9����	��A�f����d���+?#_t��fqn������g�Ʊ٬%9O$��*�u���[-L�*]� �d�H��"!b��3�C��먿zZ�ڮ �3�V׼Jţ11/?.jjD���B�z����=
�4+*rn(4Ϸ�d6�7�����K`+u���������F��&pw-3�;R�f��i�H���瘠[hb�@�q��G�&�:�_:�� 
�{��(XQ7=L��<&�m3È=UԙQ�DY(#��CZ?�ƛ��Q�I���]w��A��g]A&���_y���;"P���)�N:6쟫�$g�S�,*'��f"Ӎ���l���sԩy��̪)n�{k3�2�-���x6��B����Jn:
��k�55/�R��0@8���ۨH��/KT����>d��ցd� \�@?��n�o��V�'
x�Tg�5J�M�<N�QAw�\\�De���=�N'VM~�A梪C����a�c�@x.�##�w�9U@/}���j6�q������Q���o:�n����ϕ3Jh(TѰإ��U�C�W��n7�/�Iٽ��M-3B�(�?��O�R~,O+Q g�����ǺĪ�j.BH�/x��x	�(����k �����ez�Ż�q�Vl.���K������-f���̰�k�:�Đ���� @#q�/`(�РRL;q�ϳӚ���
�_\2�����ql�B�:	�:�d���y�G�U����H�C4����ʸ3�4��ޗ��7f���<�T���r�Qj0@�����6((����Z����h�3J�i�Uv�6c3;O�Q��ɒq�h�<!�ʿ�:�G�i��M�����u�W6:d�Y�D�:���"�)���TCkh Uf��)�"XpE0z�q,�lѓ�J� ��`�Jퟨۿ���L
 �1��w��eg���#nf���J~�H���5*G����i6"d�}B������
3U���K����6��,'7Ξ�F�������rO�����?!Ψ�N&���k�-�U6�<��h�O_W,�0~EŽeE^_{��C*i��A�`�Iw������z1G�>$wjQ
6����g���@�}p)y�{�5������k�A���{@���?����d��`��۾jf���{�A�V� `<��2^�r�Jλְcf {�v⿿?y�Qs�'x�}5�Zd��sv>�=+��uG����Z��p����� ���ì�	�s�{'I	�le$���/Dgss�"2*WO32�/���y�l*�lIX��a_o|<���I-SG�K9_���Te�l�](C�a�l���v�lآ,s	�~U�=_%� = � ���uӾ���Ռ��f�$Ѵ��#C-^��"�p0�*��X�Y<�LK6���v|r���ĸE���y�}���%�t� �a��l������0`P�d(���O��q�)o��t"�<�q:����A2 @Otl����ChG%�&���=����:���VI��}����|4���৭Swf���R�(�-�T&O%.�z��쏩�
B���� �~i��0�>����	� h����N�N��Q�&8+H*j �!Q� �^�� Ӝz�j ���\�5�rQ��'!��7A�'.C�{L=�.\������ ��K�Jw�aR*��ڍ�-�<�!S~깚<D���a��O�� �p�-�a]���g�L+�G�wq9�%���߲!z���ZX��sjX0x�A��B`$0Z���`&�R�p��e������c/̆K#���gL�m�ŇUh��\���s�ل�S/���x
h�R|�T9�9�~ݔ1k�p��D��OU�����m�A��m��e���G���w������0+�z�ߠ����O��Fr�����5w�t����\��W�D����[��@|���JU��:<{�O5��墎~Ң��~z�o-|"�@��D�z�{�@��X���u3���&1 �@���L�H]�ss������	Q�v9{Vx�f���;4qh��Xb�� 8ė��G�'QA�4Y���B\�B˱H�},*�\�?�b�v�� �ӻ���c��w�6��4���H�s7����_���s����� �x�0�Q?5t�#;����X�,p��q9/w ��$�Yp���:���7�M>?᧏�������&�mq��h���K�Lm�/;?O���-;��,��c֯R��[W�)�� �+��4 �䀦D�B�9;b���)�w���oQ�ZP_��� b-9���p:����r�Q��\z3�N����r��t9n�q�����q�@/-��J8��9��U�^G���5}tGt��i� �ϳ��&��������;k^ir�$;G�ql�^������Ա��϶��(�h�f�!'6H��� �0�o�%��/G2���r��쥓@|�8:�KVSS�Xdt8;6�.���f�M���f����#��^��{�a�������.��X�?�cz���CyrpT��>�{�K9: ���kArQz�����"2A,�|�;W@���7�`&�)�>^����9.H��d���v\l[]^V��i��@� &
-yӿS�-hי����R�'3B@?���m���kU��0&�X���h�BN�1O; ��B��"2�2/�l���z����H�O�z��0a�i2�7_3d��Ц�B�w�2�2��Zeӄ������C	E�
��^����~s�'�l"�t����F�m����$ZQ�����"�r�F�k.=��<y���Ta�|g�^�ċ��銶��q�W8�=�P ���Dk7�Ϝf��z��V���)���i�]7�O�s[�]�r X|@����D�o�	`ܤ��8�ߥ ���������n����sv@ԧ'��j	����皵��d�����{�:M��|/%�6�O�M�b������7�m���܉�%_ڟ�6��-A<u�^�v-f���Н)̲[��~�P�������#���Ωaӄn(�ڽ��%cO(��b�����w�s\�0��9)�i����[�=������	��!읃:#Rn��ƽT���$�h��K���VbJnx��4�n�9��[]x��I 翽08ts�}e��O{)�%L�#W���o�R�o�D᫏O��HG��;/�8>�J�e�1��[�h
fҤ�:��Q�6m�����y��J���N���}��2r�#�ź;)B�/�£�����U,��͏Ҭ���A�����}��Rx��P;���٬i_���.7>���qM�z�0�ۣ��6�؝�x��(�|'n�\p��+�
��| ��S�Jm����Em֎�dg�g�E*���i�v��S�tM������������TQ%`ذ^/�--�^-�0j�qSD��Ɛ��]���F�/���K{yy�p#Xg�'s�U!S�`���	����qs�W���|�c9gꕡ<pf��ڱ�<{-��|�s1�9V<u/��{��݃K�TE��e:1Ҭ3�����É�����ł�o6D�����Π�����rb�͇�-����#`�>Y*�:�����v���{����Qk:81.�G�)dI��&�������U=��!H����J*�,Ü�Z�d��U�]tGn�`�qu�K�~:^3(�iK��hy%�?Z�%�����t��8Ё��/�(���Q�*6�,�u��1�m}-r�C1��y�|�X�\��k��HK���ޭe�{��.E��B��䗛�J�5���I�`M��
�z���j��YCi������>#��
1�u�H�@k�TWjfc!d ^���2�6���]���",��#0/4��KR�	~���fӽ���dcj��%�J>$����(oz�R���$}�U ;_�r�ޛ*t#^�<�ՂLik��3���S&�E�%�:��X̼��w>ꜰ��>A��B�恛t�3�~ᠹ�I�g�`,N�	+1�B��;�i�T�C��6/9*M�`�b�OL��� �z/o�?!�)�:�q�EY��Ch���\���4���F�@*9<�x9��@�����n���ݞ��ڳ�Q�"��.�j}�- �&�>�����cPg��s2��nH���M3�~l<�������\�::�"#�*��IH��������q�WᲑl���~���"��e��ly��+�$��g�nOҖܐ��~=�q�	Mѭ¾*۳�%�\lӭ>(��-��ĸf^]*���wŦA�u�lb�1�$�U�M�"ϻB
�LHDӷ����KQ��:�8�~��R�/E���m���r��.3<�Z�w�o��~7�(��v�C�5L�=	�^i�G�HdK��,s���������w���A�"��O_`���՜ ��n��j׸���&o�>��0�%t���vUS�s1���ɆM��Ns�[Oas�Jd�8�������l;'v
e�������6�<x����α��rO|�Ǿ�}	��W/oMߪ�qB�
���)l�SE8S0@�*k�����!4��ߚ��/�
bk�>���/	�����
S~Bq+QΏ�kE,�~���x�b�f�M|!���e並}�g����uS�Fop�N��T{oT����-`A��(�"lvFnT�0�؟�w�}}K��
���h�]�̽�׎1W/;<E��Vⵖ�t۹E؄�����)�E�&f�Pg�����[��zN�~1�q�b.��"j������?SX%f7����.���N��m�W({�^ܕYgCkP/B(?�J#�3<uB���&��E�ر���̔��,�nՙ�z~��K~F[����;�Ćy@���������� �K�hBn��s��=e�{FB$���l�x������B�,�%0( d�z�I�������(��n�(�,�ƹ���[Se�V�^l�k'^|[oӵuR��8��6�1u��]���(�(�o���c5H�=E���i�k;�G�����hX(��7c�X@_���Y�($����u�#OA��[�� �����+E�n\�A�Y���{|C�'�����%���O��NLM̨��C�d>���hS��4= �X��E����gr��IU�,8�������ոK���h%	Wo�%����j��Y}5�l�ҶU��>v�7�e�.C�J#9�F���R��j�������!�8v��CW9�kW-�%� �>{�b&q��#%�I[��6�uq�e;tLj��,�����m�·N�~��=^�
4o����X�hJ��Q�6z󚝪�FxĴ�p��
,�٧��t�F{�o�.K��b�T�Z��K��l��*D9�:�K���.AdQ�w������ ��H!M�C�<Ϥ���d(��+��>�^Bn8 z�_M��n�\�t�dp��!���)��qa�8��Q�]�a]4SV{} c�9<���*�X�j�����$�tp)L믅/�����^ h
�Nɟ����C*�u�X�Ĝ���{u�
o��;��5T��[��ҏ��4V�
2j2䪑	��eF^:�~�.�?�s�x0��=��௪�Kq	�H��(;:y��h첋E؈E?E�=����Ƿτ�ƫ�.65�	����\��Ĝ�y6��6�O;M�u-��ع�K)�b��u����g��U~7Fz�[�W"��z��5��|��\���#��2�������Ї�x
��6m)�����z���Z�O���,q��g���FP��iy��%
jګ�.�My��7����b��k�/�ٗ�Z��65g��xe�t��ce޹y7�j7�p�H�^�@�TE�ի���<��@���֠:��r�V�^m7`��*j��%�_%.O ��7QU�+T]�r@�IT�A��SH�MI}7Y������LY)&�!k�,���W2Qa�U�0�ח(R�8���*M=�ч�Wȣ��NZ�<W��#�b���)]� J�����`����z3�WϠ�����]����d���x��G����*jF�6fgU$#Pd_DΛ��%��J�`��L��Dm����~�����z����b����ߜ�R��z�駋Ҥ�K����xصǼ��������ݣ�R�Fj�NWغ�r�uu^��p�=��_ٞ�7;�/�*1_�<�8<��{�0Tѩ��;Z���<�p���K�����q��r	������Ӑ^�YA�<%
���ң�I�K1�����aw�w����۝�+qPz���f�
k��i���Nj���=�)�-����(����B�{rÖ+a�p���%ቻ�&>r����U�l|��r
�y�*U����bN��T�'�bi�%Fi��Dl`����gowA~i���$��QG�͵_��r�Ʉ�2�dj��H�{��VXI�,��N�6�u-'��0����4���SXEe�X��R�m�\]sZq%����R�,?��𕙖;�[�7`R9�������h� w�L�m""}�mu��I.g��FߨhQ��rbP�����}%|a��9���H��q�c�D�U�n��M�>L����Q|���ܥ��D�vMc��#7�9�ر�Jg�ǋ�&��~����)G~�O��<�\����T���0jz���9��eӺ�s5i(H��������m�;��7Y��d���إP�8S�;9e�7O�{>�d2T�SP���{Y��>��~��c�{C3aoN��x?J�Q}�pJ#a0Y��Ļq�h���������+�3�`����T��9�݂z�{s��=��ݕ���ν:����~�S�,�Sg_�6��W��.���o�&ANL��Og�WË��YIoOlPT;ΝN�+�N������6���,���V�Uk$;l�Kc��A`&��B)f"�;��_6�s ��/�>Y01!!fb�^���T��o���r������~�kL���t��Oh2��jM�	�	��Tv��{�|C��};��U��]i�CZ��2-Y�ЊT}̴r'�>P��K�� 7Ks�3�ۻ�z�\*&o�vn���(�H�#!��+��C�ƥ���yX-�!�_�e0#���F�2-�jEg�TR>����\B�S0,3�Y�%�.jr�4�����3�/ߍ��:��Ys��s�}�H7gi������4� �^m�;ݦ�",�ư�xd�s������[�̀Rx�� l��� ��`\�n�aK��Si��N��)�V����V<���o'��v��<�l%M��!e?���)sΎ1��4�o�Dp���"k9եlɿD�bL�� X�,1�~	��/��u�;t���(�H����7��Lw.�������y���18YhTŠyA}�9��7����)�;t�!�K�$3ˉD�;���(*ݚ_q
;��6'd��Z�l�Nˉ2Y���}�i�����Z~����K�
�8Kq;�(��E~v�=���Nx
�/ߝ�����7)xރeV@���) c���S����g���iyt�)�k���PǗ��gd%����GIK+`%d;o%WD@5���N�b���7�7��Z��w\��T���O��P��f�붰��M�d%Ak׃f�Ղ�������n�b
#ʣ������&�����#� ����9V��2��/܆Z������;�#���r��F����%��-��^{Xx�1D����:$����Bl�
Mi��N��i:p��SL��?L9���S]� �40`n8}�I��ס�bz*��Г�t�q��r(r],�_��i�*nn�],������M%̓�����4���T2B5ۋy���0��Pn��xKôzK35/|�k��	58�Y��&Ll���t=�X���ae+��ث�չ�-@v�~� ��D۩S��P�/? $�/}o������p�u��+땹��D��2�h�C��zb����c����m���nn�����3��q�IF�Bc���ʽ��2>��0ެL��WY5 ���(K&��c�`������v�m0:�i�`�7_Z��������e�t��Tqp|Z8U�Ʊ�b��=٤�δC0�TCW�NFK{wL�k���zțVq���F�%�O�s�H�/���?s*�;�a�m��;-b����7�-
�>�J [6Ј�k�#ܶ@��M���T�*����x�2Zwo�y>��S)��k ��59��u߸4�Wة��.`�u�2c���p3B8�w��j������zy���/��2��j�O�I�T�/A�E�e����f)����^ d�
M��	�1	�U�����g���]|�����	Q�����8�"���������V��p��r �ma_�ի�u)
n<�U�i��>����y�ST������-OQ�ǟ�FĀ�����o�ޱ/z���*�|���,��R~=�*]%)���7��`ms;���]�hUخt]Z�p��~
ݪ��L>�S$7J ��m�.��ꧩ�?��_~}��3��Gm�LT�*�����9�m j2��3�]{�ZNɭ������p9oD���x"M�C�*�1��\��N���������Ti�R��p����')+!�O5n���#�h����:��q�!W\�0Fj��M�>(ox8�m1�>C�!|�ޕ��$i���b��k����5�jH��$S�C���\��C° �%�) ��5��S�4�R�\�IF�W3Er_	�{<������Wai�����D�q�X?��s]8g��vr��a˗jT�up���S{		+O��J��Om�6���������/;^�Yg�o�2����&�z����%���(�P[�i�4T�N�t"��5"��P��k#���յu�א��}YW�R�.Ԛk�]��V��3?6lS��ymN$�:��S���S32�)1f��ĖY�Le�|�"����$��
*���n�����Ig�3���[��L���s�(�#��1��R|Dҋ�KM�8�&��hKـ/j�P�n-;���P����@ˉOo��x��;��s���u���D���iK�|�_Z&>�n��!"U�/!Zp�̡^R������n��EGB诳~#�t�ۼ�ڞ���3
��)Ӟ'��f��y�u(�J�s�7�b�W�|uʾMx!��spl��+�ow ����D䖯�$"�@(�]�Ԫ�y�����)+��V����k��G��V��[�>�O�x~�7l�f �x���6d��ַ��Oqͦ� B�M9�A�&�F�U��V@���Smw@��uF�$�[�QE�m����d����S��3M�C@����A$�YW{-c����R�4�S������b��>EB���9g�%�;�"b ��m>^K'��B{9Sތ�r,�����d�0?)��Q�������XIp�B|} ��ޝ��t�D�bC�O.�~B6Hb8��C�&=��F^Nt.���Ꮗ�L�˻�\�=�S��ʫ_�c�����v�J���0 ��u8���s� J���;V���
�+Hx��'�/���u����a[�dr�
q8�#�$�f�C���#MB
~��:;�'�&�����A�i��pջ����C=�=���;�.A������9�z��r$u-W��Ia[2�h���x�-.�V/WYX�H!���A�@x��Q�HE"вQ0pe�~�J��-Qk Yg_�ۣ�'z��')�Dd�E�k��4�X!����o�)�����:���5��mG�H��
{1�]
�d$����{�9��Z���X����D Xm�T{2��y��$�F�䛦�JL�t�q!�r�l��!��y߯�&y,;�I���K{#��S"ױ�S񈭻10��Fw7�\�q�P3ul+k�>g����a��ѓ*j'[rmlw�.`ت�G�1�%l��6�w�#�a�Gh,G�������[)@?+~%�����c"˷�ֈ�,�j��
�7�f��s5ﬖj?�����Y	-���k;��-`0<�K�>b���N6tP�foE�ܡ/�?-���{u@���hI��p��٣j�*�Vm��S[b�4�i�����Qe��A�7��(P'y/g X���Y'D7���R��}�Q!"��I�;�����fZ��$�	9���d���NH2�&V9�˅2���V����m#�
��;��GKߛ��1�7	�}y4��J-1���K�x���?���_=��^�3�ƭ�K�K?z��!��I�F���ѕ�4�o<�:��^��4Xщ��b�W��ӄ_f�v@j��9�G�@�����l�ߺ�	������ߴ5�Ba�e�T���f�D}��ʑ�۞g���/���y��IW�Z�&1�:􍒧2�̟ӄJ_��e�gs����{�!I�x���=��a��l)jj����C��e��o�a]c�܂�����$�����j>I+��r�^�T���'~h>7WןK�Ap�S�AA����2
���+�� `��� ��i}� 'g��6@\��8}�?Z�����W{�aj���<{-`Df^:��ߗ��GI��	�q����OwcQa�%%%�G�?pk���B}����'

t�cQ��ז^म/�I�����	�X�2}��k6`i��e���l3
^Y�u���J�0j�G}��ԣe�|�轞K�Ӓ���T�[���H�kk&A>>A���'����l��m�xd��]6���D/`$]���82�Ȃ��-�_�90Q	L�,#o�1!F�		��4�r4���jjTk �B z��G�<�m�p]]~018�K#{z0�wv��b(��>*� ��3�z���D�K^�LN�u���L��%Ɠ���6���_������w��ō�������Pw�,we�M�dX%����ꞆZw�: U��c����ߍ j�6g�V
�06W8N�Ե��EQ������{�ը�z��6�._B�l����<) ��-��VV��$w��y�<=�xEY��"/wq����?�ћ���S].L�s���E�ҳLt�m�s��]���cO����DH FG�L�/�`*t�+Ͼ6ӑNf9Qa�P��2v1�E�����������un|��,�{˫K�ʦ?�(���C�=w�Oeeè+p����D�Pp�O������%����ܢu���Q\��#�h����qP��H'�I)����F�F�,�[w�:�����s亞�?Q?G���:�˝����9fy�h��n��ν�n0�+ܓ�����ɃN����l�V�_��dؽ��'��G�U�wCTB}��e��6�9ń�I�E�J����;o�c�%l���Tm��y��!u�Ն��e4��ղ���|o�=iȓΕ���QQC��Y����I�o�c�>��a܈wݳ�N�:&|n/��a���#%����P�ۂ"k���x��:/�\��|����������Gs^�)땼��[u�)j�FM�h9Z��(���|�������!i�$�i���B�˙d�Ϩ�X�X�g����_T�9�^ڒO��!�Zt�v��Ǜ6��������ݧ�V/S�Z睔
G\�F��J��9�*ԏ�Z�i�fo�Ϝ:>���F;w�u�<��a��K���c�{���T�6!���e�������\U^�G�+T�
���S	��ieͧټ�aŧ\n���W�u��'�Ss���7��SP����ω|���̩b��������lP�t��-��S��7����gf��|6Hrf��a4�/�)V�9Z�!go�Ÿ�1nf���G��-=�0��p1^��A��к��`<O	w�O������r.�MÖ��0%���=���*��Wݵ���u�̘��Sՙ��Eg�EQTQI#3c��S�VQ���UA!�C�ִ��S�,�:$J	��S�cJ)I	�s��I��y�6ϟ�~���k�����}�}�{���v�W���z���������<Y�-(�-j"~��!����R����4�s׍Ĩ%��aH��t�|�i�7��7塜?��m���a֥��9�Iڎ���]9��������v���;Hj&����Z�.mg��W�_�!�/RXt�L��'�[��k�m��ͤ��S�����"f�ػ��ɲ���o~����3 �K��������x^�W;��->��X��ן���6���ȝ_�rӄ�-I3ȅH���=Ц[p���6§ݦ����r��q���>>g��[���a%��(���j�;��qX�Ґ.�׳ܘ��̳$ڠ�s��J�ݤ⥖&ޮ�[U�'��G�_���"t3��Z[�3GFY�[s�	��#�۵����G�L���^�Ll	�V�骴�ڞ�z�:&��O�n0e�5��y=���t�+z�{X�{#<��~F��l�c&ux-U\��k��N��.�}TgC�h��� G�[5�x���r ���D3bc��4B�.�>�0�b��4H(�?�I��-��臢:H/���$�f���&�1؍F��4|��.xt
6H�����՗�](�.�#����,�y�(N�]�c箾Nd��i��U-zB����&@���*�(K���2Vs��K�z�Fٽ����֝C!w�_��m`8��E��3�ؙ�ם,��#87�)�>+�4*N�~�@�g��-�KMe�r3gֈ3����T����Ń�?[��*ئ8�ʪz[�x���z���DK|�|��ı�;�����w��q3=�R�K٥�ՑRL��I��q;Oڔ�L��6���Z.6@�k��{PjH�Hj'��s��'^�L��s��j�>s�U��Z�/�X����j{�*�6S���@6���/
�L�&2f=͡�u�M�P�E�.a'������'0� @u����s���M>�k����L����H�.���TKnEQ14ec���r"�� ��8gd�y7��ykkw���0lΙ��7��~ct[8�&,�59m4��S[�Ȁc�n��K6�-3>�ٻ�|ҋgEԣ�I���������0 ]Ac�Y�и2�c�\n��@��^ ]׀jn�W�$ϓ���Z�5��e�1����)h%��d��$�������Xo4*��k��N���N4�U�7|�H��tȗ�}���|�p,ь�~���z��;|��]����+8��		8a`�L�EQH5�:
;�`���?+^.���<�R��~���x'�=��~a`>��Y	�i-O���lPE}Vw{eV0;�j48�f��A0�l���l�k���?O?0�؝Ѳx�|�{��\��ނ�<ؙ����?���4�q��a����V�Z
���a���N$�%��Q:��~Vl�����l_8�=<�r+���U�]P�����e�c���|Fvc���v�hb������2g]��s�`�>�S�$����W�{_KcU@��fǄ����9Ƴ�jG�I��l?� �qi�X��C��Wϱ:!���V=]��7|Do�0y�|ͳ|5��HI�X8Ӱ8�=O�G����2�a�����m���������b�Hst��vIb�Ѳ�9�C��'w�'�P1�̘�R��rm�٭�<�
'DK��	>IIYY���Gh`jC	��ղVI\����H����<~Y���4��`�w�]!�t
vس�%��N=�zS�����I���e��k��hci׷�bI
���$��z�XӞ��:5̠k��G�U.UѰ�hW���۬�q3�������n���h�{��33җ�I�W)]��?���5P���)�D3�Y�a�W��@O/3K<�������s�x��j�g����6���NL��E���2�U�\��<�k Wm�q�#�>�(:�ҍ
=Shs���l8+Y3�m�ź�+͖7��NS(`�D19O3������u��Rw&���Ly�� b{َ9/R�C/ۓ��)��e����EV�^f��� y7GP�R�3�!��"��F�1�q-S�K�ǩ�����I���0`����g�e�E��ɝ_��?-FI���ŅzkD;l�f�x��D���j�!����4��`�I��L��fRX�^ї~���[x7}���-D��]�Vr컣�	mL�[Ɓq�5�V\��j�/z��#�⸁6��O�X�RS4Kp����m�|�C�5��/W֏�����fZ��v߼f��OVG�>�"�5�i`��ͷ�`s��8P�)>���VS]�*����|�y�94��Hz��w�ݐ���	M�ݍ�w�>9P�'�22�g_Z��||�	(?4n����1�A=��M��{���b_�����cBӳ�h�N�폯g?�+%��Y��G)�D��xC/�PA�e�C���	���`C<��H[K)(��H�OٜX�S{�S��~1�FW=�IƯR�E�lg JZ�0��% �+i�koL���G�</Q�0zy��5Ѵ_�b�9jf�5ð�L�o�n~�o��c�߰��z"rs]��3,�mZ:7�������Fq�M����#J�gg8k���={-e��0�C�f�Q�[�'�$_��\>H�v{��0������\���!����S��\��*��Z�S�?@:�jm�L�0 U��ȯ�{��P�t�V-�T1ڟ���Zp�l�W�(b�&Wc�����0.g��Z���dӼñ�ѽ���ʮ�F��;�=��r�T��P��Ǚ���
c1x@a��$I�+3AϏq�ځo�z��Oy�\�:��@�ژ���
 0����mG�1���"S7����x�],єA �W��3�f�a�xA�j�0yB��k�^������2�V�x�	]�����
��`�+�� _��E8��&�΄��-\��+������S$�l��d�t#�
F]�^�k��	!�X[�V&�[�PwJ�vCc��D�o5r������]P~��cd��\Ei�}��.�G�
�D�c�~A�gD�����^�X�r��~N�k0�M�KH��o��"1��iIĥ8�P��P��'\���z���Y����/�A?_�*�6jg�l����Z~���>J��0��҄{�����A��r�E
��������;u�kR�b��c�r}�8债"h3��|�դ�r��⢦�z�:����PU�6_t4q�sҫ����!LSt��+��#�Z���� �������_�;U���!T}�ϸ�2�,�R!?�0���M��<w���³T瀋�.���Ҭ�QC�6g����|��h�F�gSs3P��G��e��e���AD��e�х��%XV�tq��̑�n]���o:._�tw�X鍛ԏ��9���I_��-��#�}�Fk4��F2����m���N�p�����F�\��_���3�;�vF<$�8z�*��K�$�����?`l�\�`R�nn�t�zY�4��aN@��B�r㬵�j5ƪ,�Z�_+�a��{�s�N='�c�gE��F�mKH�sٴL�6��.�rO�pO[�D.�J����-+t]�K�χ�k[ny[�
�߷}#�+RX�C@[�Q��+%�Рy&�
2�8d��и0ʢ���k���Ȁ���k�g��=������������ D����_jIC�all,g�����t8�.M�&+j����1G�8�������- 3j���@�/;7�=s�)~N�6-�5!�)h�e�2*t��%��!pZ٬
�����/�ggo��=�x��/�k��X̴�zܐ�>���m{N�K0�RI�IaN<Q�GxB�W��r�W]sK	�3��G�#�.����oA���G�$�:-x�v�o 9��Te��rb��R�n�
�d��aQZ�ܬ�(�1�/s갼S'hޏ�.T=�g+��8���"?P�r�2$�C�[Oŭe!a�X5&���>c�ﯟ�+�/�p�;��,�?:H�$yN��a�/��T�]:�>�,���\·�'�ͩ>N��?��#c��W.�*Av-�"Zw��r-f�J+�|$���+�0Ƴ����g����� 
#��/�/���.��E���G�i��A���.8;7*ܕ�6|�[J�-:��7����y0{͒�@ >K�/7b�uC�c�d✪�w�6o��L�m�/ �~�K:��.4'i�}.���Ѻt�Vn�S5ΉY��QZ�؟��+��eT���K�+����$7���l������L��I\[@i��. �ʝ��DX�E����p�}��|;k�E͢�G��h[I�\
329��n
���BQ�u7����Y� p�t�@7cz�3Z곱���/߹ �HC�e�������g��w�y���a+ECqDckݜȈ#w8k��hv!gS��t,�v�Um 0x��i&�zt��?.��g�f��%Z�f8�� �s0���Si�3�k⁮��6�$����LQBr���+_�H�[22��6��Ƿ�YǀмЮP���ۉ/�J���7j�{�����T����_����tns��I ����Ι���P
������?�>s��Ü�H�@`m{��V��y�.�q����ݵ�OՃ؏ak��
���G.�o�>��3.jڶ�R�i���R��3'�(�q��?����06��ܭw���_w�@Z�(�Ơ�J�5�-[N��]���9����R+���Y�ݠ�q&w ��׭�q���_�🞣oӈz~��͏�!�]���2�X���n+M�VZ�O+f����m�-']��:&Dq�>�����Gf��L��N%�O�G��< �g[ ��h����) #�����E.�Pu+�*���3<|�Ku)i�����m��Q��Zv6;��{�	��o����֝@�w�F��cu�
�d6?1���WX��]��PM�M�L]�j>S�v%�(D���3v4�s�`� �Yկ ���99Buf�E��i���i���]�h
 ��i)�"Q<]�R����7�|�M�Y�;���C
�Am���zDB�1[��#���z匚�gs�������b@D��BC(K䑍��h�~~�н̝!+ ��[�fĀl����(��#[>���lq�<V��-< ��-Gq+�*&���a�Wmw���P;2?��-��� 7��e�Xg��/6ט	O
m>�����;����X��@ �y����[ ��v�^iJ�kPh�����U]<��K�08V�tm~,m+~I��f������Y:.���R����P�����f��h�WQ�S[��+ Ͷ+$8�v�S��l���%��V�%���ԝ�1!l�m�d3���ȇ�2F9嫶ߦ�5>S�y9?Il�O�%�KX�C�w�3����4x]�V D|����e�Ur���~sN�CBl�ɼt����Ʋ��t��^��B�Xƶ�)�z��K ��� ����Q/�+��S4�w��R[�����b'��,�5mb����W�^��p�A�C�eU�S^0�w�Y���;2e������\��2�6x�_����#�QY����v�����x�`Qq�.�̕��55J�=@�{{���B��'��'ߦ9��I�+ilO�I�'S%?� ��7�S>V�zU ��*��Ƌ�wt��u��$�$��g���J��}}�]�G\���Ñ���O�~Z^�"繨o��;�;C���I�2�+��@�R�8n`�N��Mſ��Ys|�2��t'��5W�M7.^�w�G��Y�eD�A��K��f�>{'�e�8�������g��ϡG~�����\�N/��	��{���v�-r���`a�y�����$k���e��z<�&������;�K;�rv�2��z��=�
�$����7�j
�C��*_�y�>�\�ӆ��$���疕z=�j���}�^ȉ�����3^�\������t^V!>�S/��0m�/�����e��LX� 03pd/]~���(���Pv�ɮ.�����|�9��S��j���]�(�J�{+ES�߀6��i4u�zw�+��^�"j�� ������:����[�:祦�E�z�6�����u���m�]�
 �y�,��Q��=�Ӗ�����R���EL��e�?l�#��{�PK   ���X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   ���X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   ���X����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   ���X��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   �X�X#&g��x hz /   images/a033a989-baef-4d73-a136-ed3ff270941b.png�w�s%n�舘�N�n��mck��m۶��m��������3��?����ɓI�If2� BAN	   II�* ��  � ,�������>8{IM'  y�X
2 ��-%*�����2^gՅ�};�]I��� xV-��H��*��rukrk��H��������cB������ن���n$�+%�F������W��H�<�:��� h�0�6�V�9 �������n�6o?�HT�1M��$BA��|�|l1b�I��*yR�����Ƅ���2�����@G��9d��ẍUH�E���ErR�;Xv����)�.Ә�;��n�����m��q�ꦴ�6_�*�q�Gm�~�F��wh �܇���A
�U}�c�8�˷����ѦG�i��#��ڋ���v�r�@tR����G���7�Y*X�Z���+y�W+����F��p�<
j� ŷ��e�vc�#�����[n��~�MB[T����ϝ��M�-�f~��=���(ق������/�gR)��{���y��F�?ɳ�O��Ϛ�c��#�J������U;<䤬�C�7��LP�I3ձ������7���>��W/����l3�,S�̅�]U��3���s��b����ǧ:��%N �mĂsna�2��FW�v�e��GD��ͯ ���V�G�HLJ�[B������60���(![���R�;u�	�� �[��̇hG�5�������5���ЫZ7��nu��^(|�-iv��ۨ�g���}ev����89�g@|��kl�=q �*�0sr��	"�6�gW� h�Q��a�����q�����ap�ܕ��^�Ϛ�<㏓�#���t/�o��\~��������M�)屮���D���ۣ�Yi��bt#Z ȍ�)��!����d�_F#$սކ��zcK#/�:!큁���u����P,��3�!��d��{�(�gcj@��Zlg,�|m�*5M��\����;����p�x�ɞ�����S�}�K*!�q�)�9C3<R�����7�s���Ľ(�F0���lx�G(r?��
�9]9������k�?��`�����j�K\�glf��v��r����$;N��B?��LаC�n�y���7��.�5"pK��io�o<��eψm�h�k\�q�):r6<DB21<���,�c������]�Kfl���)��;�W��~/h�y�������sŎc�TZe����A�q8}}�k���y$�J���
)O�\����օ�Q��0�h����R�_��{�HY,BZ�A��0r�ds,>π�)�U�,�b��^��&|0D���9Ev�_���\���*gĉ�U������h_U���p��n�#=��'00\���)W����I�L0;���O�_�!�p<�.ۤ`�C�A�_���Ϟ��=�1�A䃞��j��!���
�?t tH Ϛ$�T�pP�R�2���?�~&\��Ŧ/�Zc+�͎������@Əfz[��b �_�1t%�G�';Oπ��_�z?Xi���I+�E�S��
%4��������.����#x�0x�n�}#4��H�cA����2ݶ��J��_Łoԗ�yG�Р�J�_ۉ�R�����q����r�՘�rC���0q	cn�U�M��(ৎYD��X����녅]C<�=!AH�I*b��DxHp��	�?)������ci<�,������;X���WZK�C/e
�����D��{M�I�U���P�Y����4}18��q�9P�g�j��P���/��F�>7kR���<.H��"-o8�\��M��I����"m2`ը���&k�ױԋ̮���pd����� � �F.��|zߜtLa��Z4�v#W�������jU4&4cp.SdE�O��5A��بd��W�r��%:��7t8�Bqt	~�!���H
�o�x�{��߆�y-�b2��X�An�U�ǾV�[ ~�.����I���(�g޳�-�m�@l����P����nH��6݄��ȯ+�[|��V���xq�<��ۤy|��=��^0��ٿ��/�D����]��0�_�ʪ����N��lO�~m�1��q؎P ���doXi����w (�9�/~��ҷR��]"�"��q}?���Q#`��J�=���9��q�
�({�r,��5�{,��B��|oP.r,K{j�En;���a��Z�,��R�ӄ�QG@�T���ό�HOFo��Ԍ���ޓ<P��w�T-�,�3i��e�����;|�"ѿc ��k20Yу٨�����A�X��5l�zn�v��v�첉K�#�U�F�c��|���@��2�����,�뱷�u'O?�\����iqV���D�V7�S��cTϹq�L4�?%��=G�ŉh��gKf�7{w���-����Vd+�x{���e�c�����Q�����$��oECk6$��8w�Ֆʠ�z���W�c��>N6Ȥ��ǿ� ?���:��̥3�*/3���Y�����ݩ4{�7�QFAt~��R��Q}i,�	��"�)�YLDϛF��QH1�	���>Z�����KsdmĒU�R+$����������߀�6�ADuEa`��o��K�%��C��b1`%6 �Z|���0�i2yc��
�*�%r�,v�X��/��pH%C\aD����<���E��T�R��^���=��[��q�<PT��[I5�}��O�_g�c#����Sg��Q�`10��PUΏ�P�L���Fv߬�s�S(����!�4�1$�vVD�Ǣ���PT�T5����.$����3��gL�I�1|��?dL�y!D��r\��ðλ������
�O�İqoPH�Cy��:�H@�(���|��k`e���������m0f�Vݥ�Q���S"Jlr@�\OWA�ȏ�Z�$}/��T��gA��4{j�'�>���.-��]ye�{ҝ�����"%����;�CGz�'�4{Z���Hh?*��� ���7
��8 \�g�y���Ja8pI�!tqz�f�[Z�9pU�rʐ��w�e(3L����eю!I����`�ظ3+}���Q�w#$�c��{L�q~(������4s��Q�{�:ڸ�᪵s"�+%:�Ts@&W-�5�{�������5�*�vޟ�@7h�7��,{tq��3�_��1�����k�"i���� X��\
1�_eedb� �	�� �|����n�"?�,�*:���!;XS����(�px�6zC^TM1\Gy�
v�Z��c�
޼���p\T>�ڗ�K����3��덍���G�����Q���s���A:���Q!s�7㑱'q�t����/q��X�c�"��0�0Ö��2����v׷��ͤ��j���&��ct�.��=�=$���s�T)����h�be����3��	'>�}:Tsyau���pcc�C���t1�i��er�=�~�#���.f�yL��! f��X-�54p���� ^��],�/y���$�{W�G��Do�T�h(��Y(I��)`�{d�mٓ�����}�Y;fӉ2~v8���������[J�WNA����i1�>%�'�yMAu���noip�&Q��9��.j�5��>[����9�3.3��Ǎ�Z�	2��ԗ! 忶`M���p�&�E��M1I�����+<6�: s� �g�VjK�Ԥ�_4�o��:�E7�p�(i,jmM�V�K�w�0��H-�L3��U�D�����@z�9��T��ˌq���M�Ъ���$�c��ދ%�܂Y���*��J�AQ��x��G�M�����}�
8m��56�x��l�D��<aEV���C�®��DW�yR�v���GVg�RP����]�\N�of 3`� �>I��g8HF�m���Ė�vV�}�;g�-|���1� ���Sˋ5T�K�ʓ�R��Jv���M������v �]��;�	�#~����#.��o�!�aH�]�����R� ��>zXM$����^����q�{��r�6�y�z�oP�S9Ѱ����辟#m�R��źP��flswe.�?~K-�vgM�:h(�0H�,@�H����Y�:��Ͼ)>��b�#�M3&�#A&�%�R��?��]%��[��0`m 	�H(@���ɇ {���|xE݉@d� ��
�|�q�ǎ��,���@���Z����F�0���1U�0��ɍ��caveL�� B��>ĵ��|�|8]Y�YbF�
���:*plO�֡I����T�m�,jk�;tU�QxΌe�~�M�TO���8�ٽšU3�`�u��]4D��!��'J����.�t�{�9!� #�pc(=VCS����&7'/�Ъ����j���f�g��� �t�a�4�"�2�3���}���n��ܮnNmbϜ��|��+^�{-�GN�`��.ױ��U��ʨ���a�ʦ[.Ɍ�ұ���PT��ɏ�cG���@�F�^P,'U�r�l���L����FS�]}u��֏ӑ�_F%dc`��[AOb�_C��t�K�|y�Xv��e#vL��?�����;Y�Q�����(.Qeo�D-r�p�����B�a�r������)O��������H΢S0w��l#l������#���X'$ɴW�a������*���%{1C�O���z+��H]=q���
�
�,D]������C�4���5�H�,D>v�x3�[�t��)��#2F�_�%y��6�*e����^ts$G���~��SP��#_�\8��Gb��� ��FR2.��)�3��8ߙ�p쒋�4�w��}Ek�x��H�|H��%I�Ĥ�I���C/L�0�����k�N�2 X�c ��x�͘�Ӻ`�yq�= `78�p�߱�Ĭ�D�����gLB�K��D_�(,P�W#D�.
b��V��w(�_K��Yßgp�ʸo%F����dn�}�R�G� �~��eXԓ�lj�Z<�R�l�gN\Ԯ�̡���/������E*L�*������LfS�	g��e_
��jZ���)lr}��� >��0!��x��̰�G�	��Pڋ�tō��Bʩ?b`I�WW��qj��oE�^ܬ��Tfظ��\,�����7J����4b�H�	�) (��
�;P��Z�L�}`�!���I�.������E�4�L����'�9���\j����*��6��;�x��=P�2:9�3F�2���m+:a��9�$FLg��M{4E���x�ې2�?[6��{��n��h�"�r���"�I
3]��A��U�)E�.L�b��M��S-G���?��"0R�6���RyFx��9�L����H��\�k�0��=>��^߷x�ܵ�k9�%��;�;}s�>?"z_��������y)��)�"H�|�häf_�Z��e��b�a�/��N2w���4iik�H�^��'Ҝ>Gt8Ԏ,;c�D���=�8>.Yj~�Tɰ��x��Żz)ךN4!�w�r��Q��a�����m���P���!q��#�W��k���Ш�����T���
|�d��R!�@���2�n�I�rq��`�q��8��@�L?3w��49�2\ֻ(SJFQ���)����ˇ�]��t�*0�(r�:Y����{G[�H���4�G�!�����mW�;���,�%�TJ­EI�`���g&���0�!���/�ЍC��\��2�d��e��5�evŻ$R`JMtc���^sGp�f����nb�JaP�=�7�y�W�Ф>2V�)��ݻ�Esg��x�eafT�rE�����Q��ng���7gE�[�y3cM�-�lřњw�
�WE���R��s�n�k�k���� �WR��Ǳ�ߵ�W�h��!9�?:�]� ���tYך�k�)&�tVb��[5�MM�4=`2D��(-��}��k��ew:%�b-�$ބN��2X���fʐ|!��76��rb�}��� �{rNT�JMJ��wL�f�3��8E[c��Ldp�����؄�)�!�'D|�6��T��6"�0�j�+DS��XJ'X
5���zVɿ�qeš��UN���.�k�Bh�=���	u b��a���F,�1�O��	f��<eD#|�e��C�%��1�Zh�TȻ?E��*AwP6��?D��)~��b�m�aƪ�9���զ�FޡCk�u��[QR�%|$Z�12���?�%��D�~�lo��.�^�M֎��K,w2��W<�E�][ ��߅��^;zN��U��!�D���'��A���[�,�ؤ������_zT<ϧBt��������J�*�E&:�8H9�@4F'���+#ԕ���4l��l����^4�ݸ���vڨ��n)���\�~e5��	t�͂9�Hb9�*PWH�<�����*�������x���z���a��\��a};�c�]�?�A��BЊ���ڿ;�EX)\PWi��O���|���ٵZ/�3��,S>	GQ�z!��
i����3����7��]��=JV�HW��a2�O�?�QB�Zq9�
�J����K��ǂ�C�S�Ǘ]��*��}���*��Q�x���1 �a�	���h��Z��8G�P���U�v�<�VS4G�^�۵��%V�7���ܗ(EV�����^L/<��-I���u�r��Sa#������;?���*�q����+x$R4=�!Q2W
��"�����1�p�[>{��'����/�&����G�a�����R�Ht@��:����I���7��*iX�U�</`Z���>ξ����k1H����Qw�)s0�CZ�S9�}\9��;����1{_�P-g��,�y�)� -��_Bv�_^F���d2̉��1���ͅ�!�� `	�S�"\�;�O�C3Ķ�3sT���AjR��K �e,I��O��Tz��U���d�����d�O�k�k���x����C�#	zO��d�+�Üe���H҉�W�Z0?�-Mm�[+3L��r��uO=������<_NXWU� v���qq�^�T*�N��hI�!�ؠ�t�p�~�^�N��9	�J�1�b�9�����
&&������Ĕv�F��J�7���+ZM�}�*1=����,^�.0>�l�bT^ߺ���i7�fe�b �y(#�GEI��`�@�~]Q��4ƿC�e{��"�3�'���� }��=n�赘�,OY��2�>:�9�Zӹ�8\�X$�ǒM��D"��pfL��#��ߡvU���
%7IN>�� �����dD
7�Ƽ9�\4A���ףr�i�&�rg���6"�f9�>��c:�_|��YX�g�S{�SNQq,��hF*9�^Fv������T�� j8�Ee�F�y�<�t�\�Xl��$���{ɋek�ku2�h��$<�_����Kʂ~��Ue�M߼�:���D������O�r���L$a9>#�����$;!�`��89ErL���}���Ah�r}u���Q��;^��r����Ucz,/�zL�ńG_%12M�pI�HF��.j�V>?���po��^����V��88h2�o����oT�L��k�U�xr9���o\D�#��>�hO�~�dp��\ ����+��4CQ�~&?��]A# CǮeɝ� =�8�	V�Xe䂏r�����)0�.�*3D��>l�}�*���p ���fu�f~�}��p�K����J��d�r}�@�hՔ��תo[�:�^��V[�!��p9�.w;C�y�l����J3���8^5�g���� ��Z���	�WM������g�oRv�s��5�����N�|����KN�R�Ł��n;�U�q��Yqb�"#M���ͯ�q���2oXb��"��?2�H9�Yul1�lm���ʑ��
�t���5ߑ��h��5"�2��g8y�>x"LV�sa]��l�6�)���s]�d���9�����=pP#��g�/��e5�p����y(���+=ޭL䨼3�*2X�[�B+���y��7�cGC�)��b�3[@C�8�m�� i��S�Yᨄ�I�sHWX�
�Xˁd7�آ���ڽ�z���	�.%M����d��z���~nשҖ�˟���t��:�D��F��\����t=�Ú�6� =��`Z�X���i/#N��R���K�x�m����i>�F��q���sF� �A��W*��ֲ�r�f�ǘy�O�_��ȝ�!�@�X�i{�\�YW7S�ոPP��4�'�����kh���0�gC�B��]N��Zۂ� 4�'<�����d��5�1O�J "H�k_p���B����~y�э�+���R�D��sD��iWꙔY6܍�N���T��s�6l2�(����H����m[��e��S���2rsSG��W��3'Zm����H�9�q�#ud9��n�dtW��4���w@v�"r�|vR.2����#'F�I�b+��% 5j,�L�Sp���*�d&�4���m�N���]l��g�x�*�g|�v%�n��с�r�4�4s���bzQe�m��>1��z��4�>0;�4��ɿ��p�v	�S^\\4,���
���Y-62c5Ȑ��ۂ��y�mj�34𑷔+T0����r��{��MP�ӟ��]kYcL��t<Uv��n�-&��{![O�d��)pu��ir{5o[��r[���w+��� �ÚW
R�W�Ǥ��B�<Ԩ]]B��n���Z��gI�q�o��T�8�xa_�<P�r7�K؎Rī�:��.�Z�~"
Ϸ���&	3[Zf������_!������$#����Pƙ�i�F��F��G�:�5�(dy����Њ�ŧZ��L��_vJJ�hd�|�!qlV�D�de�1ߩ"��Y�0�lt�1�Z�v�P����,�V���v�X�[�I������&�ɭ=�~���x��\�{*p��ݖ����[v:IU���u�h��y��v��%��P:C�J�(����R&�(m�L�d,����TB�>����3��n����G�I)�>F��S���GLF�����-�g�9 2*$q���GA�����5CMl2��B_@.�6�?��A���r;5�#C����K�bj������7��M�?x�n�e�������ef�3��$�MCh���nG>���?���1�n� �\�>���crw�~�?;�!��9���D+��������{�}�!
d{Y��A��
D�d����SA���ˍ_�5:�\d�]Oo� ����S��B�t,D�w$o��Y�e�%���Wk�,�����Oz�.J"� Z ��ԄMX�o0h�իnn�,F�"!�c�R�#%�,#�	}��0�����n����Į��I��I]�-�0;���0�ӱ�M�dw��xl~e8�E�Ю���́�;�׈�Pc���Ż�g�D"_�+�]ߌ���
�:�Vd�	w�q�#�0�%.`"O�F@���D��	�����B�N�# mv�x��!T���| k��ֱ�������gIm��s�E�7���j�� ӢBkFă���}B�a�IOyHk����x?D؃'$טE�Lh�Th��LA�'���k�I�]����qR�zT�{n����f�.x��OȔ���'�7�CU�Qd��0��V'�7����������D�h��/�Gˌ�<u�
o8�1H%r^��Pr;5i5S���L=⦚�q��9{��{��?�ϡ�Yb�iv�;�W�qnOϝi5�E#�Y����~�2����)L��`����g�`�K��|b�8�Z��M�P���������~nԎ���]���jE�a���.�m�9:���s9'˼y,7 ���`�{�>|�K�>>�+ؐ��H���	2wTp��5��ݍ�d��e �!,���BkPi�5���I,��L���T����vy����_;��z���>���b��$[!˖|zIԀPBA�#�{��"T��-�F�(��H�^�eU��YT��5j�y|�ʌS'����+�ce����k�j�tU��A�3ƞ��rY�������@�~��6�!��.L��+�Ǻ�ԓ�Sm(\d���������dt��1{i��`3
�r"�;�
#Q6�/��R�˚θI��M$S��8X,O��k\�'��z۾�H��r�%�����딸Xh�^r��Scb������֌��>l=����'�uT��Ef�W�w���6�M���>�>��x�⶝�ޮ�˞֋&�h��Ҭ��{{��<��>�ܒy9�~矵
���>�B�xPV8�	���n�tW �4���ˊ�,���y�0��@�1M�s�	l0�%�2GDE��h�*����S�y)�W\e�	��܃_�`y�BŢr#z\�_,ƨ�b=����PGv��a��F��5t����:kJM�����u��'�p
97.�V�A�w}>m�#���e�mT_H��&�����(7&P:�a-z��(�	[Mѽ>����>W��xa�6X@\Q�h�lVrV-����&��e�_q�
�)+cry�ry=u����]�r�b�RG�����,��H�%���5�9�vwC+���("N�����7}�z��c5M�y-�b�L^
*4^�1�u1=��� е�8,� ">���?���������u5��pu(m)��t6R%.�������JNX�H��7�1�M�	ʖ�(򮖄�Oޏxg0��=, �����}�z�W�x�c S澽2�����V��o�����C��zڗ�
��+|vCf{+���p�
��M	'�iW��S�ǃ�@t����r��4��C.�?,�PZ�d�R�+����%��tG�<��� �]��̶�L�E�_R~�zp?4��{_�&t��dv��p��F	�t���L,-�zn�q�.��q���0m>���*��q�T�z̟�=��%L������]YHS��.���$���O��K�b5��(Z4��L��#𫕀�V��կdf��*N�v��u��}h���ۼ��X���h�n#�������ѩ��qI�z���&�A�)˚��(73-J����e��Y�
��TF��ཇp��Z��qt�~�������^���u�Õ]9���M��lz|п뿱�Y�y��\O�"`/��8��G���T�^ݵ�]��ѿ!p�/�}���{�m��N�؆���B�e9A�g�j[�<Ѯ�w��d�@I�o���	���=�Ia��s�SI��j�����ϵ��{Z�O��m��9���������pU]��:X�~�GY�����Jf���Zؕ�
�`��w�zͨ�-O�,�|��2����yNP(ta,�u�F�9�����ˤ�sԚ�5be�Ť@�M1<|��E��R}эf	����UO�#�����85���y���l�M���i^=_	ʿBX�5=���p��s����n�����}NVF��4��0��O�H
��Ɵ����	���#j_'TX����&���Xd|n�L�Y�����{�<����(J���w���?�(���k���ֽG��տ�k�[�`���'�,n����5��z�5�p��h�/�K$�;�>Bnh�е�=��2��ޟ�Ms�*)�2���壱D�<�p���{��
8*��}�q\�B�Z�ND�����
D����W�!�X 
���>R�6�=2�>�l�f����}G��9��Gx�B�/��j�8�,�uݙE�\<�P8��^�:��'{�'����'��l�W��Xr��R���v�fX��YS��]�ʏnayYՏ_��Q�	�lי�9]y���dR��b��$b���\ޭ����������[=ڔ81��_M=0��$��Y�_��L-�C��� W��������B���N�=��O�ΞU����UD��x2��T��HB�'U�r/�B��CN��M�������6���y1�������ي�|M���c�+�}[��,w�y��]o�_�[��8Hj!�U)ϑ�~�Nc������F�aծs�,W|p��/��c������`-C41�����@���L
ɰ����xx���#���,�U�$�z��A�`W�u��J��{����lf���2y;�B�x|�x�l6&��q�@�oK���cmwBChgUL�}�&�&t�N�-��Cs7����es�R�ɗ*Fݷ��	���*��ճ�h����c8�dI;��~�=*���Ǡ)�%h���]��S��z�d�p���-����.d�Ev��-��q�b�*
�7���;E��R}�@O7^\D���}�;���$/������F�0�zǮ���
�g�}Yf�@ ��$�����u|;�z]��F�Y�ھ���v��V�$<���"���,��l�ν��&�C���r�g����T�hd�*�z���+o�#d��y!U'(����	� �eF���䗽�r��k.������ ���ſ�^���u?���{��[�Z�{�A�J2OF�4��¡���ʪ���$��&�ne�}�TX�ee���L�v���w��n�[]�����,E�;L�쁿�MH�hR|����QI��ẗ���bΙW��@^qŧ�-��!t��1�b�4�蕿��R�Q���:�>J�ƜZ�
y��f�+v�CY1x/�Z�-َ7������Q?~	�J�"(��QC�ڴ���ՎØ�j`�%��0�ř9�l��&�M_g8z�lt�fC�<�J�į��帜<Q���q�v{�ؑh0	22jƚS��典�@�%��}�<|kn7O|�#N`��vj�{?�;S��Av�k�~@��7�C�����vt�����^C�+����ֱ��l�=��;R��%uт�2��{���%��|�6�T�:T[�!�=S�G_^vi��G�i����F��������Z*AC�<*R\��~X�*���� � PU�M/t�s��p�W�s�f�DOCW�w���/���%� �t}S!�o��!�������x�7���{��͏���DD ]�+Kႄ��}*�k�6�����(d iRM]����ȱ^�(��yz�t��x�)�g�rI��eK$�ݰ����h@> �$�k��B��� ���|/O������X�	<�f��[q����D�(�_��^�mIf�?��|E�W�{���G|�W9 %(����ڸ�X�ā8��-��'z�+�옌����;b U�y� 
+:+j��+��}�q��i�o|�o�JQ5��J�XË�]�/C�6O1!}����l�_���'/��n� #+�Ʊ��{뺋���#�����Z�ύ�{�b�9�:�ˌ���c�ҥ����8�oG�W�+�|���K�4�p��%_x@�:t������r���<v��F�.�{^6��I���ïN�G��+���tfj`H�U�-�1�Z7^�n��F�N�	�F�u�*O�]U�8&]z�߁+�v���#x�1#�����%��tH����ၘ�:�Xa����f�7�@��`4�+^^"8BX�sN��D�����8��i]O�	W��*�I����i�+G%�����?`+�X����:��ţM��'S�EC
n$�`�=^�]K�������c�����B��~�(?���fBʹɳ�~��!��ud[)� ��!���2�F_���T�vw�m�{����N�-݁d�֟#�|t�3��,,N^�n
����$��o�G�w��z�y�'^.is�`�0���5��˥�V��e���Ep�׮��̬w�|謼��Dӷ�M�Sͨ�¥N�v� ��r��*ɟ������g_.4�0	+�2ԍ��̈�"�z�����=�$��Ƀa(����](�Bvat9㢈�x�K��J	���۱ݜ쟑��7���q�M\L�@���M+G��=�b�o]f�zOQ�,M"�)�ps�ӏȐ���+�N^����>{�P�nV	7����q�ִ���$e��EdU�x�][F��+���o�ar޷'W\��D��kם�e��<��q��B�/��J�����E�E��^��d�Q�B�$_L)Gcu�}�9�ӡ$,��̍����s����ͭC��"Fl�SW[e���<^�=m�,ld�i�<"�K�p�a�k+�)�J
(�l�!�;�eRf��uxP��	c��iCj��!�� Kf�]a`D>cT������X���F�n{M�.�vA5����{���M��b��f\�*"_�o����Õ��/�r�F!��bd�CzF���D�O?��a�����ُUZ�ͧ����G�h�U�nmݚfv�b��L�ʓ�6�N"�1C��Iw�2A�j͠�#o�t�v���a}S�^�צ�0+�FJ2�]i/�DLY@$~�)laЩa4�ȄaQ:���ſL��t�<kF��)t�-' T��1=�t�!�P���&��Ӎ6�.�{���X��5��cg�J)��@V{:�
p�@-pe�$hZ��)gH���D9ih��a �}y3;mdP�[˘].���9����(݂�o��S����G�)�.O1S3�B0b9��}�@}�c������=���:Gf�ŹU8z��G�d�	TD����G�j~����-�qӭ|�j�Jݐ���$-��;�9^&ri�1�q���h�k�NK��[��Az��
ѯ��	åZ��	���-^�-��x��)nh��Qux	ٟ�C���%���8^��N�,���y�8�������R���{�u�2E�,#n��wR����d�(A���[�ml��|��7Y��4БaIc5�$��n�u�OvT��)��(8_�%�T��D5ݒ��b�+����it��I�\S�e��Xv�;M$S��`���>��t�pm�	AT	�����n��4�t߶��Rg^B��\ӡ���h�+�!��0�=U��.@c$آ9?�z�`X��I���7.��!��Y�L���҃]gS�F���DhvO�q\{���6�y0�ts�e�Yh�/����>�*�����T���g\�'��[��}��1�~���]����@0b�J`l�8]m5J���S��>F�e('���Y�b��&..��%�L��Z�|�s%�w��,m��,h�j�6ׇ���Jz�E���"ZB�S��ݜ��e�]�GS�2�N���ėϣN��w鼏� �/���q���o�-��Ke;ǧ�ú���ӷ!)�K;-�ҘR�0�ŏ1V$���hg�&�iY7��2��+�]��̟]v&���G]�g��XԢ��p���5�Fpy~�B��=�{�p��б���0���_>>�f�h����.z���q���U;N����Ր��^;��&��
���n�u��R�������eA6zo�.EA�w��47J�fYK�4�����"P�e�r`�\=j.u��B���:�abSE�i|�`�d߽�I���n�Y��R�Z@l:�����z� ��RY��a��ʋ��E��ȴ��j��!*ۯ�l@����T,]T%E�� ��������i��u� �]r��@�p������r��\_�{��_�S<�d6p
�=bd�)x�� -%K��C���s�"�"��_
>�3�c���� `M���"7�M� ��M2���Q`�>��Ax�� �;~ĥ��7 '�9�-rG�'SE�)��^�����)��x|��Ҷ�u���)��?t{'V)�IM@��II�n���UY�LL(�j8!}��^�!��ɕN�<�������m��F�8s�#�۔��N�����,Ȏ�U�b~s�����:5�y�<@���f̀/�-�Y���?�?Vn��s�k��dM�fH��ڭ�&m[���l$b��ퟱ�&;XE'�.�xC�:aT0�Y)��}LVܛ�!.$dzT�y�,���F},K��g��B'̘x��|Mz"�-;���<pi��r��n�x�w��F�K�'s&ʿ�R���d�_�o��P���&��o��=E��r:��F}�����7������>��2�e@���| 	qMW��
W��?�S��ħ5��=��.�}̲�9>���w>�'����D��UB���Ci�����e���{J���^�P��u�t �L��l�,*���" 2�h�4�Ax�EM��������Jde ؘ��aEY���=-5J�`Y�_���VR��Eb3�L}��c��pK�U\���;���(�7\W�Ԗ�X���v�%' �Q�i�䑝0�o:�aM7�th��È<��j���1�STc���&X�F˱Y�=��L B�� @��Tn��"�A`<	�	���	apE`̾m۟.WW��v������?��?r���{\8�����har:�9#VE/z�El�Y���)�/p�n��l�-,�Ӟ�iK��9���M���wm7�#���o��γR����BAZeDaR��T,6f���z�^��������~|��uS����}�R�n�p���c)憹�Q�"�+#'��w�߮왭C��.���������<�������ӥ���f�
p�{]�{1�l�� L���HR9ma,�yDAb
�77��g^we4�����R�i¨�X
���dĜ��Czc�s
���f����)&FA
��ۡKEO��<{ʾZr~*r��G��v��hk���f�'[������	�ښd}�0�e`�$G�cUW����>9{���윒�x��u���rUݖ���ֶ�C�Y�!���r��Cr��cx��ƈs���A}�suY�=�i���<���X��g غ���!��Y�]|�#g��Oaa���B��i��_#E�J�%Ҏ�ܮ�kt+�r�A3=�$m�ǈ!�#� ���R��a^���cnF��zf�Y�JS�Eօ��E���1�� �5���Lzԉ�zf�q�c�qF�\_�{�ԏ�� ._yrafNPsc|9��0{D����}�{q������=Z7��-/oꍚ�U�����> ���f�܆]*,��)`�n=�Y�NȌ����K��$� ���)/mBgGܱc��"����o�p=�;�Zf7&�,�+v�f��s�a�3�T y^�9���$.���)̛����Du�m坓�?*2�g֣PS�tRk���mT+�
�uߔ�P#Pt_�~u1>��zeN뻖�,�� h��o�O��.�1�3mw�2��'�\�~]l��B1o:�B4 ����:�<����g:M ����ic�U&z2vi�Z�(Ȝ�?�Rrw�=�G�/�W�"�� �тZ(q*N���ۍ��߄���m���7�IN�b'J��2���ߒ�v#�_9����&^�������z��_]�{��zթ���)�.<;�&� ��mͿ����v�A�Q�$m�EP`"/!<܊� �ַ�%�` �
�GyH��^E�_��3�-��{��ɓ����}'ٿ��cC�1���8��q����)���q��n�}�sr��y��T�-��]ݮ�y0]6������w��u+���������//�k��s��91i)���@�>0D�Ϊ�v=��ݔN�cC���O��0�����S!tr���n���U�~�u����:
t���O"���Q1Ff�����G�<A�9��=PHU� �{� 2F8��Q����%�.���g�y�G(�*w���L^ժ�\��g�vzV�.�B��!g/^�1�ÿ%���,:�^e��<U�{��Q	dk�)�!a��(ƚ6=��1��.\�>=B\�e��5��������7��\�!�3Sj�lm�>]+k��Ʀ9�m�5Ke�~��p�tc�`[h�!��0�#	��U�!3բ~�ͩ7JE�����l���FjnfFiJ�)%�Up� �~�Ϧʔz�ӲP��h���6a����i@�0]��R- $�q���Z��pW��"�bE=�}���_YH��ۈ�	��Ņ��q�uw�#���!��k�SDl'�Z_�>��X���j�1W{�ԙ��Z;�^?�a��h�vĭ�� E�����kFX�;g��"���\״��̴F̧�gts�2x�έ��W��5��$cz�9u��x��a�3>�z-:6�s�nQWt����M;s3b��C9;� ]x��2\_\\��n�rR-@�S/<��ʹ����y�`N���SÁ'� 7��#q��f��:�lcZTb�o��
�5m�0U�~R���<מ�j��q�1Y,��M�`nV� |][_�
��*�}����:"X���+6 ���Ac^�,����@��c��=��Μ�K��k�Da��^�����x@�E��#��{~A�����5�B>��H�f��F}�@:*�b$r�6�h ����O����k�;1�2���CM{�x��8К-���|���E��k��mH��~}$eG~HtkR?��{��=���u���4DN��|�ؤ[�8�n�̨�ق�q��ܩ���̇H��9L+'7g,�"��̃Ǡ �B����FQ�˧��+�z*��8��U��dK�2:�6��ܟ�We�/Ǒ���ck;���� ��yr�I��h
k�__6B�q��y���;OȻ���}�`�sg��{Uj�i=#LOЬVf��k`3��y��{��D��҇��o~Ks�4˫��n븦S�S�t�ǖ��1�>��Yw�pˊ�����~���� ��0ʳV�q����9|R����;�$7R629��D�&��HwX��
��}����Cڴ��t_�Q%H��F��c���X�qpK+�Y�[�kBor�V�a����eF\�v/��Z&�=S�I�cP𝝒�6��N�A��	�t�54�醪��T٬,��z���;������+ԡ܍���ڒ��t;5w����m��:3UԜ{s�-Gߦ��E��W�p�j�)Cfr�+h����.6[Zi�*բ�^�(ߒy��GzXe�ʓ�����)�6Pփ�0�Î�[�Qy=w0Q��<���<��q�v��˺z�#��2%�lQ�a�8�J�Q+)��uM�)�<;&����]����f���w6׵�F��Aƍƛ)<���J���S���%R���nM�0�?�����2��an���~x���ԫf:����U�3�oa@�qcEw�0T���(��E�`���>�'�Sq���sj,��R��!I��[���&Y݂n )�r����l�[Pǣ�<��ǥ0���%9����G$��*�͐g��OGf�<��p~�^��h��X��1��zE�;q<c�ή,_:��]<q��󰠖�]�s .�	 8+���E�C'��M��&�����M�e��U-4��1��H ��F`�d�0c�q�l����h	f��'S �����9Y]]�5 �!d��5��}80E�ܺo'��V�Q4�r��D>���r�]���勺�g��.y��9��xh8N��Q�e�|��ь��4�-��ZM,'�<&W�^�:��X�U6�-�N�(�G�>�
 +SY]o��TXH;�:twM#���~� �Y�x�;zP�~��פ�ik����)����	�f7����n��rh�n9r`�>tP{(ё�l_�zEmk撜ѵ�M�"+I�4T�yD϶��2Ж-?$�%@�biq׮w����>�E��Ϯ���:��s��o�'����Z,���Y��Mu=j�䁵��>�^
���C�,=��|n�֜�M�Қ*"6����~zz'����� �2�"���6͜9�)���A[,�;�='����΄�<ɾlD��˯�kl���?x��f�+��PL� 1�����Ǧ��F�૬�)�\Z����W�}������ihe�j	�U� �wM5`|��K�3�I�y�c?��Y���ԥ/������=�U�y>?�O�V�G�!a�(_wS�p5s8@z`]h���3J� b��et�����۽s\g�T.LO6�[����6�
�Pn�����	�PG +Ӳ���G���c�����5�=����&xmc� Owe�N�,���Q��y&,Į��Ls�oM��x�����g��̞��P�"��Jki}�;��6ޱ} 3x�3U9rd/[�'����q�>y���������d�{�a�̭�	���u+3��ic_��g�9�o�h��x��ں��*k�R�Xf�?�в�w���Cd��1 �T=�c�߁9,�׺�t��~ok��R+j�d���DS�<��E	2�̓�A���+ {~��N�ʯ_���fW|��E����W��}�x�%@@҃�=�n���E5���vP�f�҃��]���,qF���FyV�% �>���N���_����;�� �4��x��}�3r��Z1�c���>0�@�\<�@k<��4Ԣͱ���}>=r@���4b������&�7�'�1���B�8��0���td���H��]�!�䣋�demC� u����l�@���}��d4�tb��ge׮M�p��Y��ؒkK˚��2�f��de`�����ƺ>�z�e:(��������3��<;� W�]�z@���{ñn�%��ko�Pf�������X��t�|�&�z�qu�_�.���F�[ǜ���KIj0��ޓ��:�`�ɧ	��#�c���Mz�>�X���/��FϺ�F�E�]u:�Z�9��d������Fz���^_��}�c��O=�����;�ѥ�۽��yn��<V�y��1b���P2�;Y��&�������3��=/�[��pFu"����yT䩙zM����a�B�KC76�:#���U��u�f��p#�p�j���zF��h<o2����Q%`V;v������B��tK�JZ��&V5�0�)�B�s;/�� m`6J{��rO?%x�s���Ȁ��YZ���\��y*�SR!��g�>z;��8����q���h�������*\��"궺@#0<�UADZk��dl< b3�wqݣP�ﳘ��8�Q��g��[��(#>��#rǝ�I�فm�e7@�SSl[�B�|9�򳥹9����˧�)�W�������.-x�O~�G��{L�<�菀�ʫo�F\���a��ޕ�@q+����s���/�/�)<	����ɶb����D�&}Tn�{RD�^��lq$H�a]���zDЗF����p�4�2g_��p��:�@��/�5�E�F��4�~�=����ޯ�Pѐ���tFrF��M-6�r�J�hJ����p��m��$���i���O�]\�+>��]����7N��Ŏ���fAOw��tk.�k��E5&l�6�E2pp��;���3�\�S7S0h�Y`�������G����Y7F��ܵoN�'�v���@>=0�X�h��~L8VOɣ�-��C6=c�P��R9��W��n�g퇭ug����Ֆ�'�0��dO-Vd�1F����>�R�}�`�7�oa̖WW�s�\5��x�'��`���!<P����	��x=�戵|�Y8l�ǎ��xV=��F��b�f��2W�Qbi�p�� o~A�ɢv��ck��iW:`���w{}���p;���N<)���oX�ú��U��؆�w �o[�����c:�̩���n��-���׌�Ӌe���9ִk`6"0�9�in���Ece]��%֖pV��t���.���Yt�����6�Ә3���$��Lk}U�0���� m4��c���
֛��8����"��zSS&�H3�]uLݳ��$�s��c���|��1�m(��e=��P]k��QcE��|�.qkH����>�D�i�H#�t�~cZ�N��M+�Ӂb���ʊ\���;�(Wt�X��b'^n$��Rډ�?�P[�Sձ������_Q��{u��s>�M�;�Y�����6�$&k�Cx-�/��l<w��n2L{�E��Xt7e�d����L9� 0���5�rL2*v�8q���?����T��1[H�Vc�x��ݮt �,�2=0�f^,$�M�CC"N����R�c�L�WNx�VC멦���
�5"��M���5Jb�K�A�f�2w.�o	=Q�&����7���J��2Gn�6����a;g2�)�K! 8}��7�!��>)�������Py_���t J�V;���0�fj�anN��ե�,ml�Օ�lB��	�_e^6�m��˧�����wJE�'�zcQ�g�E��R]=E�p�!=�V�̕�>�-�f�bd��;J��n��&R���Dz4 �eN���>�G;�&&�7��Cf V�ou�VV��Ȉ�*Ls�oM�@�����40������0U2JV��i��ȧg1`i�H^��+��ҕ%�t�v��7zjH}`�����C��a󦪆t�%O�%U�3Pb�llA�U�a�l-�lu�2�n6�PH#��j�m�)4���Y�˝�j����5Ym����q����3pW�m`��l���α@Z0p{��FZ��a�u�5 �����kb{9���Z�h�&ͱ(��榦_fg�4Zr���ZSu��%Ϳs��E�ۺ��)4�U.���Mڸ�%���6ܜ��g�0˟}�~��9��lm�1����v_6�c�<Fl�0��NIw*��㵥됻d}eY�(�W���2�}X�����7��U�,�Z2���Wʳ�m7��M�v���3�P�4��]�|�tU-W4���2M�㴙���gZډTO��vzz�b��N��&n�kM���{M��-����-�溞����^�­�0�<P�ݫ1�h�Ab38�d���y��k����G��;s�=y�7�#�i(��x5*i;ڇ�;�(S���X\���o(�˱������̲�nz��EP�� 	d��&���t7{f�3����	�D(b��~H��]I;i���ӎl��	Z�l$A����ʪʪJo��9��"��"$MoG��1 ��̗�}�wϽ��svl%�g���\�|Ψ��3Em�v�~(�+�A�#H�0� �?�G��l�m"�U�^�����L����� `t�.��������1� 8�	 \�f3ٜ|�ɧr��e��	�9e)
�e6i��GZM��?P��Ia�Uq�)@�z�PI�~���dhhH
����Z�ڙ4����z6m�$��I�}G�c�B�`���[�;�+1*��
R��Ť;����0y0�y�!�Y��8;;�:��:�����S�<�5����X��}�Y����>�����p�lWc>�M���T�KVS�'��zUT��[˷u����/.�� ��Y�`��؊�%�O 
'z<��ƆE��3p�ˉ��㵽A��̦,q�&�h��'Jv��1�'�`�N�t�\�-��<�ԛ@ُ��/��:P��6e�$a:�J31�R�����i��!+�G&B]���pomo��W�eF��!�_e���@����K2��I"j���'��JV��ݏ���K�H���������g��z^z�z���
9�.�������g_r���lU��w�������A8���eת��*��E�6j���M
�����f 0]�����`�7bˀv�0���H��I��/�X6��|$�+h��}}}�f�i�����F�s���p��1= �4S���ẩ�+�-9ȩ2�ʠ��0���1p}��u���P#^GAƦ���'�1�#��E�(���?��؊�e�;�Y�u67�Ɲz׵Pez�}zA^y�8��(zX6�E]#�9S�[�:l�8rcM9�}�Ң�7�������^VI����YX��Be �/I�`mp�p���G5A�guM���4���_�xIΝ=�l�O ��^���U����~wCפ��R��M�DD]���ordH��l���=��Ϩ�7�0��}D櫿�%��}��#* �664���؆�~��ia��& p!�SͰ)  ��1�r� �_��,����A�tj���q���DE��m�d:GSR��!����&��e��#!ҭ�P���HV��F�����:�~I�8*e���ǥ6d �~UJ�٫T#�Y������Է�h��.��5i�kh�閵�2��#h��Lk���gY��#PI Շ��(���Y|��$1�@T�m�253SL>!�O��~྾m��%�.�5Ԋ_�YbaN�0�����f�F��.�Z7��]��)'~�k��3��ԭ��E@]���CX��������q�{z,���g�
�ib�|�Z8�8`j��*"���p,Q�ܢ�GA��4LLϰ-Y�˺p�l۶��&��Ρ�/I� xO�?&�㤠|n�:,FU�Ƚ��ҡ?ߨ �T��yTE�91�ke��/!���}+k�W�� �_��-�"��5�i�b������,�*�^�[!B��VV٩���*�|��:�nE��f=�0ߏ��ܯٍ�i�@�,k�'FEM[ɳd$H�� ̅��,�<h� ��%�ː��C��{�b�T�:]F.����R�tO�2{waĀ&8�ZF�| e�\[\	>6	t��t��+|[�4��~T$qx"�����*�|z6�)8�/J�ß�奌7��5��j��l��P�	���#\CG����z/� Y�8=��^�ɿ#�f�pB����U���o�L.LUk@�������bI6�*�n�t|A��(�
�Q�"]n.��K	#��6�-����~P��*�Y�ˬcz�4j,��X��Y�)�:Z�?�'(�����YY�����11�Q�l��Y�_VSz �:D<���l�0��c����$4u�c����փo�Մ�J\ô�54I��/��%��:(~���@����?����\�s%��l���!c�,A���e[H�5�D*C!-�=����6E]K�L�/������._���yQ�е��l>�V�Z*k*	e�����x?��;�O��k���oi���g���!���+��#� �W�h���r4x��=��vP��Q �=�?��3S\/�V2E���e���y��;��tu9����.��C#�ȃɅs�eX��RlE���D�.�鶷��E���(�;���!(]Ts
�ڛ���^&�Ɠ+�"�o�I6���! �ON�`=� ��8Cp&�'g��1�p�PG	�E���u*+��1����)]K�$�l���L6�u�$���d^3�*2�U&_��K�
���-C�G�
����i���u��(��T�TB�����Z��³G���E��=��.iRfQ�C����E�&�x��L�P �%��|��O=Ǔxz/��3���کf9}��R}�F�5�C�� ��5]# �U5����x� �������P$�*Z��t��(�W�1�H�S�,i�@5^�����<���r:�ۉu:��9<�M��ϱR��"﷗`����8+4k���s�ETRV��֗Dm�ёa���	��eX<SxaAR"��s�N��.����X�u�
������P���-28t���p}�C%I>ڢH\��X�߅�&��ze��-�;�s@���}��2+}��������)������Ê���q��Z098\�5m�Z��>��ţ� !%��ぬbppPFF��������<��Ȫ軠4�/Z�Y%�!>4�r*H�ְ���ƿY$o����4G5A����Q0S�K[G�ԣ4�Yo�f�u�m������|3&&@��aQD�Nk\.6;{�����A�HT=`q͚��0XAc|�(�p!����I]\N�,�D�	���iN>=��!aT��<�̈́�㉝���*��t|�t�
Ŷx"���|����������[�Q`q;7�J�+�?�� ����*�9�? �_6 ���@�aȵ �9]��/!�S.���q��#P�l:Ñɼ���T^��!=�Kr���z�<U��L{i}��#U�Jld����@��i;�bA���i ���p�ư8-��d�U	8%��L͍+C���)�Y3NTĪ"ռ.?�O<͒�)�7����`oԙ���
�!dMo�m$h�య��"k����v�''ߣ�'Gd��0�Ȃ3�<�<
�b�v�t G�\�Dj��y�@�|���##$4���t�4�s�Rk��)��Ѥc9�$��I������+�H���/�>z_��կ��;	�Zu�MN����Q@�̓�	��7b�-L��5k�{�s�nj6���?��r\��@���$T��nV����PI�I���+A���r�ҡ�����eyi��^gPj4���!f&JK������\����VS�T��6�C���1��
���h''��0�_^�UT]���gRV�����d(���뼬�4��Íڭ���)k�t�,��;Z)1}#���Ү�V�����h�4�#zή�3}q=c�5�cࠡ��u���@��&e^�m�����M�޻I�_'itE�i��]�K�� �'�LVG�dey��U���5���'յ�28|CN��D�k�4bI��/)����=���ƅ�t��<�k%q��i٪�g.~��
]z�@��!'�0����κ:��Ex��Y��_s+�Y"�h�m�
9I��r��5�����ls��\p--F�ɲ�7������Wl����	PuE�Xŵm۶M��_����{��8������[���%�a
��kI_�^�g�"�1���3����,�L�޵+����������@���H��c� 9 Sb��������㴜��9<���@b*�X�W����#u�=$�rL�$Ȃ-<e��xzL���)����m��,��ھ��L *h� � C��@�	�����2�r+�3���s9c���޺��FЂs3������rTH�$4Jl 2t����$�4|�*.б�)E�e�d#k�衞+��a.k�_4�绖Lʚ��M6Xv������(M��^N>����ý����)���{K�����=��2
��1;}��x�����`�M�c?���ƚ��㷭d�����H��$�[�h(J��L�+�T<q����$]l��� ������p�E	�1k�1bB-@����0��QB5j���e|m"-�q8��՟��t���@czf�m%|�$&����
<� ��HѪ E�B���7uHcM'Ė�p�Ҡ�}U"81�2|N���,�D^l�\��9L�M�����;�� ��9�A]����O��VYX����z��T�E�bm=�L�<�-�<l1E���-�A���&i�=�R�_#�X��[���ˮ/�AYowy�	�iYנR�k������FZ\�t�*��l\!��\���� �Ѥ��&���z�7Iu�Xuݟ;����4���5Nʪ��f]�)��D�į���<{<W�%�����D��-�}��oiP駹��-���&�^`I��h5�?��qBdlܹդ�?�`��V�g��T[�iF����zr���s?F��O��{�]�IL�Α��$��9#����M�.B&>N�js��.����Bb��K�<Z�	Y��2g��d�e����;=E�� �%XE���L�
���+�g�8=��"�@��sgfz^�8sQ3{�M�B~�)�]^�A%[gd� � W���I��ttS^����W��.Z���I�z��W��%�>ۼ���Y��z}P����@��Y.��o�ɡ$q8�p���IwW'�I��E
�a�=�K�.�|	VT�gA:���겜>�)+@�����BnH�q��؂��!�A�Q,��&[O�3(��9Y-+�;y��#�1���E�.ښA4V I�_A&�Uxx�aU��U9�އ�@Qأk-Rj�V�?�I�\�Ķ�CcL�"�q�
�6N!��-�3�~��5�I"�WպF#��@�`��5�.�V����[��6�K��^L�[cUP�p(B�D+w]_3��C3qGJ��92��a��Z�M�%1���]�`� A �Zl�N�&S��i1�+@�3�_�� )���R���J�_N�P����p�����+Yh�,ik�7��+�H�[&n��+��1��r}�����G�Z��8��	c:��0��X*�:v�sG�c����מX��*���3�_#`�5���=��0�ZXZi��ybuxOWu���58���Nl��w:��� �2ֲ�U���#0 ��&���\��3�^���IѿC �0���a):db��
Ø ���"�y����AE��~��|C�^�4IШx`�# �����%G�T���S7*H^CX<>$a7�a@n+:��219Jku��A���J�%�����b��d��ƀ�Ӡ Q-h��Q"kh���1Dr{dW��=8��.�Ygh�xm5g)��3�Ό�Z3f��/\8�q�����˱e=��$��4�㺮W�����)�xg$�WɈ��\-���ᖡ7X��{��B?��˙�++[(`���Y_�a�%���ԡ����,��ȍ���y���z)������&؀���SU�����Ÿ6�S�8����'Z���to���N3�� ��3�5����;��:5x�3���
����>��
�x�YA+����ĸD4hF|+Y � ѯ�M%DM$=H���`� �?gm�R��k<���{�rټ�5�8T����:z�����&��Q�hT��Һ��0��3A�¥ˬR������ ?��@?�����M>C��;���_O�������,sR�!LKR�4�(U��W����g��xԟw�����>�4XD$��v�"�Ycx�ʴ�R�o�١JZ8w��;M¢߇�R���g,�F��83�^.���)@�A����Ö��nơ�T�^E���sS� %�T��]�G�>J(�F	�T�@0���I6�F:�i|��Ɛ��� g�k't>7���o��Ė���Fb���}���"�OA��_��5��\��Jطh�g`4�J���@_s�F*C�J/�9��m&p9Q-���׭�Rt��s+�l1Y^͖\i��BW@x *b��*�j����e�-3�HGJO�|��m���A��)��΍�S��kl���y���'���`�����8^ٮ������PEN�c�e�
"ٍSAF,��1o.@I�n��û����!.\��{�[aM�&k��S���P)X'���2|rʘt�!m���Y.0�`�/�YtW��|����o�8������X����W�.]�jaqe��-o��cnNtr��N3^� Q�b�d�<I��3��P��_ ���N�n����3ȑ����& V�+��������DD��.
fܖW�fdy}����uG�S�uV�UA3BA��a>�]L��H
�Zs:r,3�V!�WbY?�(��N��\�>�G����e������SU5Q���4n�z�D�؜}�8UK�8���s��s�V�X����*�M�M��ǴO:b�\"�'�L+[�dU0ۜ����P�2+�7��h��MU��V����$��l��;TWa7���(��>���"�ԑ �D�-	<ߵ���Q�U��p�Λ��2uB�#�%�'�T�=.C\���5�����}�f�����[�X{)����;��Aɾ�����(��4�!���t�]��p�J肱aV,I�Є
��yS22�hini�4��Ĥl�Ԡee��0
j@��c:��Ѐ)��z0�P�S4N��3�!I����}S6�^@��ٵ{7�!'?�T�V��J���4��C�sal�O��~��`�aLZS0�I?����Mt=H�4Q�6i*�b��<��� ��*��UM�j@�oo�N�ϭҲ�릾�(��Ӏ�t�N^�ٺ��?L�b������5=���^i�쒚�����A;h�Z��E=���7���'*���"�-@�E���֬Mp� �<�#6p�حς�u'��<t�Vo�w��!�]�����w���Su�u����^���#}�7�7�) �.�ZXԵ_���t�\���I?���G����h���t�@�.�����bO������H�331&ը�"�ƞ��̳�]�_���D��x��/\rBYC�F#E�cx��]��n�������כjZV��Ǡ��6S� 2,��f�P��
*�Q�r���f���tXt,u03,Qk�� ��^�a����T��+~`�Xe�*�x����� ���[�@V� |T
%c�[6�d��.N�mʖ��(�~��ua��/���\�!��Ud	��P�ؑC�"���'nz���y�+˿{t�����������x�������hD;
��`�A%��}��"x�dKn{�G�*á�9�T9~�v�c�z@���@��f�X����>\8B�)! T=�E�,��\@���L�׋�܄���Yy���eM�����{��H>��c�np#`à��d������!���P`R+c�C�����Z�?�\6<T�0�[��p���=�u���nTv��)7��+5��}[���W��v��!O��<M>��������wm]�}�������*w�y���7dk�W^��4#h"� �@;r��_s�Ӭ��A3����q������_~�~fw�41��N�qG8�� �5�" ���E�9I�Ar&k�{�z=pw��%cc3�$hb�*E�����`Pjg`g�Ѡ�j�lh'B�e�ޛd��]�j�������9�<3��^}!��8Qc�<�Qf�^�K�Z�([�m����2�:z�1����/IsC�,����-��z]#V	�r���aA��
[4ZM��={�lA_�7��\�]^��3k�&��]��|qV�;�`"��g�P������xh@�z2�+[��N�R��ʱ;� Xnlj�?����[o�8������UQ���e���ʪ��&&s�����]
�:,^]W�
"
�QAL+���<Tlpq>a����4�B�h0���ν{d|j�&x�������� _A��b��M�Be	�7p�X����Z� �&"{�ܤ���\lY=&-�200@0-(�"�(�S�ࢶ���)��mr��4�g�f9t��݁��2�)N�'��8�h[k']��f���Yߧ���J�EA�b�~{����ڀw�s��߰�Z�� !���t=�eya��$�w<B�q"����y���g��D���[$\S����T�8�36H�ϒ�h�p�8����HFԣ529W����٠rc�T��X���&W�~#@�,>]�R���%pV|n�e/2N?A
6/�r#��҆n	�XL�8]������No�< �ˋ)�"Dٍ
��0�	6��/�\� ��E��^H�+j��l!�D�7��'E< ..�*��8�.��
\l�8M��j�bY9̬?���F�k�Xf|��3 =n�`��oit[�6�+�tlܠ+i�<+F�jʌ 5�
�����#L���ڦ�ɹ�_z��ŗ?~���[�?��?�z��㏞��i˳ɫ�E��9Q�������&��D�M��C�z$nn(�"�����4�"�<��#:xL�@����b3�	3�*�˹���sWG�z��P/H��Y���)y��侇���a�Gf��<�(!���nIA*�bPe��Pe���7���� d:p3�$!p����.[w!���Qj}~�P����K(��)����%���^��z`�����+ _�ɎmI͒B�*r��"Bo����T�rҩY/�\�}�=f��=�M9v��24�O�"T?p�a<k�
�]��c��t���J|��$�kW����%����?�;͸ur�bT>���6~�:eU��q�(Guk�kX1���w�V��; O�����vTz�i�6�W����,�c�7�ղ�����I�ޑ�?��,��ߓ���}=L�p�^�R��*J��>Ŗ֤��K�����R�� W�ɿ����@�9z�v6���I�P�ܢH�G0T���A��@��9�f)� ���sg)_Ϊ29OEr��LK�R����<GF���M�zTAe�kVU����9P���Q+lVV�O��0SG�_��8s^y�u
%>�;ߖ(X�	�Ug���;e%�D�8C����-i G�9�j*
._�3g��Lwʎ]�F�g&���")m�5���8)���K�+����'��Z	��9������K�>��?�<�>*���[�z|Y��
��ئ�Æ%����Z1HH�Q/uZ2
d�x��LN�*P�_��|H�8Ls�Z]O�o�l�քt���M��b�4h�����g��ǏˁÇ��M�z�'�F�>=_�f�l�I\E��&���G: �~�����=��u�B&^ �"������>�Zh����k�Y�)@��>�q}�.�g���G�}
� 0'.� @�F%:��}KR�N?���X���j�G�d)��$���0u���e����~k`�7T�t�ZYdv�� � ��S5(���;3��ˢ�ikp|�X���Ȇ�52@X�ß��(9M%^T<XBq�6�b9�I�'}��A���'@�ހ�=ÆD?��bu���0��*RͶ�6��@�X\��w���?�NQ�Y�ihs������ �D�X�D��i�ZE=���˞�M����D��Ҽ�Ō��)�,�����	-�s���uacr�AV���jF3�����7f���?y.��>��O��vl�@�#���9���+�?z�g�ǧ+9�[KN�/��E%#�WA�h�؛���)�f��E�^h���o�e�!�Y�V�p�2�](0C��:�� ���j�~���\bY��[��ؓ�f�-���p�oߵC�l�B� #�`�����@��X]é��a��A��{'	&P�衇��o�)g�_`����&b��S _��-���<�:(�444 'N�G��Ν�e��| ���n�n�������އ�ܪ�U{[�>��x�ãr��5�vmD���3�����\���y:x�������~F��w�ڦ�h53P�F�����r��G2:6)/_�M=�������6@ ���Cn;z����S'Ya�-�Ç*H���.��'?�a}���)9i@?��T��*J4蓃w�c�>,�վ��{����	��n�ݛM� ci�o�#9���䊍M����;P��r1���{��;n��2�)w����ay��%�@etbZR
dG)�����:Z'a�t��A\�3==��o?ũ$�DP5�}={�\�p�c՘�A�4�AeV�&��Hk�1����6�VS&gTD�N~�)�Q�Q�}CG�LS��]m4ČC:^�m�+��f Iuu݌�àpE#F��h�85����AbcK\�ݝ]���*�m��>��\�>$�P�mMT��N�5�/�I��0���\jU_�!�<p�l���4��ϡ��#GU���_G��>]O�2����zq����[��B��N��%?	�.+h뀿����=\��1��(�tM�5��䍷ޗS��|<��h�Fm��%�<|��w4Ы���N��gȿ%���kba���SJ �o��&��q.a �_�1o��ə1�m���	x�P�����Vx>�s�����Ye �E�V�E 箶&yR�G��-2�{�ߡ�@����j Ӣ-qHT��U���˧� �܅�^��{v�-7���E�iO�NML����JL_��� +.e$�]��4��8��
���P���l��id�1��-����,�c&z#�e��)5!ʔ��6��h Xb &�����s�� ��e��	 aAO����������B�d)���E�I<Dc�W6��M�j�H�{��q�g �S��0�%!(����pUPp}��r�l�SX���@ 4�u���9K����=��V�QZu�K)SՌ�7���d�����	�,�2�R!BuF񄜹rq��h<��t�����������{�:�l��4-|��p�'g.����<�Oֲ�;2%O�~_^;�3@M���ؤNVK���C�#F�ղ'Ir\Y�)/�"Բ���@5ePV��^V4&�Ga4�vFMuT6un���ߢ�TuU �f��ͼgh���� :}�3�r�/V�68�����"�~xTK��K�֑b�k�����%Yprb�2�8�F�FY�'��e�Q �EE@	���L�H��z�<��=̐^�%�<D�2��չ�g��ŋz�dk�.ٲ�[҉��[B���\�(j��.i�^+�kI���z��S�z?8<��.\���{��=yTv��Vd�����1r{{��/��x��UId�rMx<��h	�p ,��%9��	V �>���7�g.��{}��IId�����F��N�@?�RZ��+w�y�	��kW��W_P;P�y��G���ǧi��R������'?�}H�7S%Y����h7��σ�R� �� �OO|����pD�zu�,.'%���J��ڕ~J�Gnٶ�[�k4Ý���1��vv������ޚ�lьx;0�� ���� \O>��% ��[d��\Bv6.�+)}��r�]���O1%)�~ͼq�~z漼��	\[`M�y�d�?|���" �T?����9z����m峽18D���0#�8o����@��8� #�৮Z�T)#=ݍ�?5����iMސb���������w�ׇ�S�>���q������s+����D0����-��E!�K
(>?wI�uT
��ҋyNNA�U���JX��-�efv�{�.�ua��Kv��F_��7H�ݪ� @ Xl��Q��i���^t��*plnj%�҅s��f�(�B���� �..sﮧP�hr����*����Y	3�;Ѧij��Ox$0�)��]b�c�.�[X߰��zҵG}2�I�������ep�_�=��j�sgW7��鳍����ϰ
��T�9#�³���,;ʅ�3�����o���K��<��)@�! ���9L%D,���A�?��}Qf����	�^fD�Y��A��n�"["�%T�L�d��,*�øf�/B�8�>7Ge9e�&����&r�ʆ�0�\;�"�h�8�e1H^��Ѳ0dK�ސAc��i�fKE�C�g��I��#������w@�u��E�� ��E�/4~ԃ�H��Ǘ%��o���0�7��䊣�v�Wb՟]��?<z��>��?���_�h��᛭
��k�rS�I=�bޑ�T����g�_^Mޡ�gw��nF�.HZ㰀�QN��P�Mn�O�VWW��<���H���q��"a�:n�큲(�~ѶY�,v6���{�X8���\%Ny�'z;���O>$��Q ��k�����t�4ȃw�F6ʦ �z�ɯ^zIAN��! �ab��6K�T��/�Ӯ]{䛏?����_�6���+�7��*�Sc��ݮ���;h-�S=���S`�V�]\# �!�C3�!�D,f"(����ٳk��a�i��6ڈM�����/�ԩ�4+��w�!��~��ٳGF'�9}U���dM��t��jji �I�B�_��G����\���^��g?���w�-����ꋚ}�J,f�ccC{�P�4T���+�h���U]_��#�<����v�dAc:���Yq�űj��j�	�L�$7L:�y*�n�֧�,�|���ٙ�e���o9"�w�����
�����~�(H��tXn>pH���ĉ���o�����~G9��9�@���+�YT�W[[�	��1����L�+]�m��,͘����ea~Y��nٵ� �>P�vp:�I�j�}�~�'NPI]Sn��Y�} X,���'�<��N�GZCz
8@d�鳈)X�%*]�"�������w�4�v�ԟ�v�Ǣ=���`#鐧����N�~�Q��x|M�Q�}�3�o--����J&�{��������ʗ`/Q��d�	z�y\�x^��^��2���Ĭ\��V�_�`|�	+=�ђ�H0I�+�˸��>���Qy��G�����A}c�h�'A�ճ@�/��@²�R���^�%4C
��Q����_���_��-��_�ٿ����)��HF�'H��-�7hO<���Aޢ����騲tnꖆ�fNw]�xY����jB��c<���X� .N�
�� ��D��6�Ƨ��̹�<�[:�v+ʺ8�
(B�&R]'.}��D���yӃ&I����WS��i!��`2
���JKk;��kE��d������s����/$����;r.��_��OY����R�ށ1Ђ�$�����gi�	���XL@i�����
�Y���@ /��)�*1��ޘ(p�"lz�]�nϔͤ��TP�Kщ)�23,�ء��W��iﰠn�Tb@.�ߐeZX�9џI���6�\�Q]��	 ��e���|�G��� ʳ���^_����&z�hey4{Fpu����x�Q���b��q_0���d����ާ@M4SH�I��{c닷���9J���5���p���L��v�#Ѽ�h����3X��;R�-:��4B�
�Q��-�m>b��Ef����e&��Y�&st�V�Ľ(�k����m4o�ނ�_�J^3��fm�vn����C�M,��7�ȶ�-�'�_����� ���,�j��#�?��l�i���1�k�}s7�x���5�����a�)�˯�J�#zx��AX��gh$�˧evn�m�=��}�m�N�ݣ���}p�������  �k9|�����h��>r����J\�ٱm'uAj������������OeyyF8���z=���!*V�P0��]�@���٧��󗤣}��z���u��)'[NʩO��ɉ1}�I��n8�?��M/M�}��5��P*x����ޛ���
`�]t��3����G��g��{��� ��g0 ��$8ݮ���X�~��W��>m�J-�f)v�ɡ�g�~�߿��gJ�z��\�V��(��a@��֊��Vq�M���0�1��Z|�<K�H�$V������R��鎲�Zj}��;��D
��<�uWO''F6m��jĵ|$�:��QɈ�Y:�&��q�h��>��� �9|^�kgUT��UDe��$���7�|[�
Ы�.�ҳu/u�&��58�XU@�)���^ü�&v����χ�����9&�?� GY�>�����C�� �l�M@	�p�v�c��'U��UV�a�Y7%���6����d�����c|�������B�/bx� OPz���0 p�^�?����z
3�+�����q(�:��E�Wvq���f�pT^���s�)8�뙸*�
4A\Y_K�f��=K[{�<��Sr��[�����*�´b��P�>R� 7*�olh��H���l}��t]b�A��wu���Yưd>�3g�5|�;+!�q�8[t�),����:�;���|��L�p�J��_��و'�,Ꚛ%�@œʋ�铴�e]3�J�F��7�聕�����x4�k@)iR.Z��F:�#zl�R���lا�K+-!d�ȼ=w-
 ����%�U ������0 N���O|dq(�9m�c�~Q���r����;�H�"my�3bfם��а��w���I���/����^��<|����5LK��ύ�߆�kƤ+����e y�S�oN�Uzm���	�w ��И��E��+`<�$�2�Y�R��u��fө����3��gB�e�|�Bm�/�׌Ɓ�$�;�4=3�!d�%۩��+�#�P�Mh6�IH̘�q�m5W��V߆�ϗnʕ��<v�DAn� Q@����[�D��r�5�����w�w����AK͆4s�ʬf��n�\B�jò2�{��)w�}/�a�S��������L��ImC�f(Պ�Kr}���+i�D|I�>�aU�����6)����������[�oߦ����/�KWW���?�,y?~\n��&���Ҋ�&�ʂ��>9���Ξ?'��z��ܾ�
�Œ�?@�~in�փ�1ٺm�`֒�!�tiv� F`k�YM�'W����|��!$�Dm)� ��+�ܯQ��}�qy��(����s��jdjz���Х�4���	YX\f�Y� �g����!y���Xb_�֭�pI�P��a��KRf�p�t��&=<pր���Ȋe��'�XA�Z��#H��B!ݸ+{�.T����/dώ>9vh�l��s=�2������K$�$�C��G�t�`T5P�� ��>'W���7�U��Z�Ihh�����-M����/a�cS��7s��T���?^��k5cN�V�Ĉ�ŧ�(.�<�TT8.��l����J߮}���'�Ͽ,Kq�&U+�J)0s����m�ݖ��;�[5��������w����k����%�����Nȥ�C��<�njF��A�E2�?씕آ�V����2�^v����Y�Ț/$�>~�D�������K��i)b�@*���3^����5c?���c�G��HU�ֲ���s�ʣO<%�������k\��TvؚU�w�9�e�h�+�	�2�{�U�ʽw�?��?���:I*8���2����tӟ�W�
��C��"�mL��(��_��{������&�|�I��_>�[5�+IZ����P뤭�0Y�3F�  ��/|T�kr�ɪP�ZP|F�YR��)D�t�xp�������2��wH1��/�����- ��c�	#�������y0 ���8�b-��Rٙ-�o��7TQ�#�5S�2�8�hv��<d8�۶�jH� :���V�9n�q-ր��o��&K_���}0�J}���N�L�8,��pAn�i|a g�2V.���}L@���*��@��W���2.v�UT��� 5Ma�_NpU���~�$̗ccZ>C8�*��a�����H�[�r�i��� 
���s�-�3v��lNI�6�ϠMf��(���D��'���s8I
��%����Y�o�C�ҍ����4 ��j����.�1�sP3�5o�ulJT�ئ�h�`�Mj�� �*��W@�� 5�>�A�86��h�aT3�@��--M��{����^�f�������[z6�'�������}���������|�;ߖ�#���褺����ӏ�?��g���,[D5(��?�/���w �NOQ���x1�Q������;8���.�W��l��g����W�Ϳ�{�_����|�{�?��������ʱY�J��4��wk �P��^�"�5޾}��U��1�X�	�=	S5ܙ!�VV�-�4y$~�ZVb��m��Z��q�L�`�y4��G��'���=!?��/dvqNB�a���f�<��i��!�"�#KQ`��0�H}�ȼ�N���P�6��8T�_~�]X�@��bw�`�`d��:(>G藔'��Iq�ŕ8K��Q]��6A�+�Ϥ����y.E^xf��$q"��z)���+���s/���aioj��鑎�N�ol�k�f�Г��zKz�)R�~�i],��v�P� {TWKˌ/>;�@�e�ni��#��}r����P�v�t�0����Gw=��:�l�"h�-cRȀ�4-`�q?�*����t2N���{w�3�yZ��)���\�}�U�Y���ZR�D}~�a���(�^d�Y����.��i�)�WV���Iں��5I�o�AF�4�vIA�XI�e�1%���(�[WС��>LR��}�~���<�k�S���?��ҷ}mGJ7��.G�`�I7�$*K@�PR������^rpP���X�q���Ġ��ǆ��)ZK6�K�3�(&Ѷ����� Lz��v�m�M�=�������e��=��	���_��;A�C�<4�9��&�F�A
@2Fu��;�%�+�{�G�+��#��լr�~�AQ<e[`cҴE(� D?7�#�p�8��z�6����rP��˵��0������ ~x;A/( 3�G�=~8Q����$��S�2��ݜ�p������_q�G��ĀZ���UQ��e��*�n�'>J�g4�b_��nCতז	Xe(�zH�W�pu�L
3p��a��\eLj��5a�� ��c��?��Ô�66.����r�/J�.A�@����#�+.�m���6���3���瑶���}�ە�/��l6OǞ��򯿬�����Q=0�0��-o+�V��r1R�e�p�tۦ{���tM.�Q!B�(�/�* m���,j5����M�	|�:���0�D�8�����P��bW�̸4����"�ʰ�r���*��/�G�7�����N�{,3	f٤�0ׄ&s`#���:��W%���bRSdXK�F���;�I�LȌZ��Y�{��j���IMc=?gX���=}���/�WФY���������0M��l5�ȯ�p���Vf�~�;�<@�'��|d|��<���eu����:f��W�k��X�����D`��p���V@���A*D/{��>��\�rN�ݿ�Kimk�g��}�{`�l޶]��/�b<�!�'�'�@����N�����'�ܫ��{�����;o��c��X>9��>c͞CQ	@ O�J6e�^���D�?� ��JµQn.��A�@����[+��֤���$i'ᵽE<��y�����wNР�g\G40#5�Fo�_�?WK0\��Sm�~]�������iAp���sR����m����G����'?����jy�w���D���N�Jϣ��%R��E:Ֆ-cXҵ��\[dŦ��G�_�^�!���@�@I��v��e�4�u0�M�*$);�:v�IE1�� ߻�&u�p�8/G��Xb'$y����y����-�c��)��{ߕ��Z����ˋ/�.�U}�>�P�4V�7X�㐀��9(9���/��1���7�~G.]��I`�U��n�-����a�5F�u�x��Y�r�D�
�:�����sr��r��iẆ��W�U��2���O]�l.˩0�6�g����>:uZ���}|z6�����رY�>��I	U�r��([�6����y�sg7|�ju���w��H�%/�����C���C��O��5����^y���OP�����!�/_�P�E�s�ჲ{�vV�s�LO�H�F�5w��țo�L2��|���=��k
8R�_-F+��c��c��+k����T0w�N=�Ђ�����.㒅�	*n���7 �L�9<l��� ��X���*��Qin퐩�)�{MR��B��/\#�儔 r��b��+O�a�1��E]Rn�MK_�e��R9��l�P���CC�T�i�2��$�9�j�Sb̊-��(#�n��F�FEA�Z!e;8k@�Q��(iZ�!�B�m�q�
����P��K hTnI�(�+�� g�5 �b.�~�_7�Y	�M\�p�`�Rp9�>����hY0�$L��B���uU�g4��A�*n���k%бɼ�S[N��␍ת����$�� ��w˔���ɱ�Yb�P��;GC(WMTSʅ%_#&�ᣛ-��<���꠺�i%}�hj
D��	�*m �FX.p�YyAu��0��R������,�@M���e3�^Z����=ҽ���J�fŅ�G>��#���79������sB���l=�H���C�|�s��,���]���V�d�,M�]<T�'e~aQ�f�m@�3���3��PA�r�+k ��l�\���0��Bwm�f��l���a?K�1��c9y��:|��k�773+�h��7�Ian�&b�
������}�\��O������[HCk#��j�`j���ƪ\(�2��4x�x\AI׾I��}7�L����L�L�@���t4��~�;ҷ�� 4��"}��d�ҧ?� ���3f5;������&"w�}�^K���>����Tl�bzw�u��v���S �Y�Y�y��Q����T^[k���w@�_��?(�=��f��&�jbfA��+���?�g3K���n͒�%_gp�G����
�!}.d��kZ��o�Çɧ'?��#+{��D?��,.��]�nK
Pܩ��͐�_�{	a8����i9th�4vl�G������2�(28:)(�#�}H���\����V����q�����u�KgvZv�O��"I�.�<��!��[�����'�;|!?����Q �4���a&|8g�TA�Bjط�_����*R���{e%a\�t�y���0TN���I0iԹ��ܙ���u_�[O}[6u���/� �ccҷu��n]�"Kq:'s%�-�L��3� ��78[p�N'�edr�� (</�����Ss���`�b�V��\WxR9K��@�zG��u��tv���#�Ҫ�br|H�[�$RT@4+�s���!�ܷU~��P�r�T��PG�ɱ��e��A$�SҮ��Q��n٬k7%�Yy���%��������
T`u�sQ�����vSf�G{�v�ҷE�{4x~� ���g�+��)�$���3��1�.E{��i��Xb|�t�=�ط8�En�&c_\��d�gP�g�Ŗ@>YH�]6�+��XU���^�N_���X�`9������V4�� �E&%|t48����{��e{���g�*]�$Z��aO���R�6A;��s��r�V�����$��%�����Ԇ�F�X�-�����3FB�R͈���fIt�eX�_Q�/�:HK�A�/,K���J�@� "� _�8ŵq�*S1���l��d*fT�m~�
�d�3�
X`Fh���Őo/�g  z�X�mm0l�*�h����r�ꢇI�C��Q������&��:*�䔋��ZT�g���t{�_�R�_�����O�6�f�;*���23g�3ZӨ��f����2�t�$X� ������20x]���w�����������d=]���?�g�ɂ��q���(�N���� �����M��g��d	Ft�L��勳dtlV3W� ���6�s���Hf��q9�<����/����
{���ă2��e�����Y�@t���{�'?����xQz�o��{eێH!c(�.���O�h�t��=S0�50�D�բ'�xR3�ZѳV�%�.ȹsW�����E�#�֞=7ˮ]7k�ƔG��N.��^*�Y�FF�����������S��o=.���S pL�}63;���"w����9{EcؿN�a�v��#r�}ǀ1��=ăvxxJ�G'�����{���;��Z�/��^�g�k���A�t��lgJU$*�lJ����tv�c�"���=��bY��}F^{�]ʍ��~�����v��:@��lH3�&W~��������F���&phXY+�ɏO���;���*$���
w9�	?���]���<�M�g�9�'�*� ȖK�^h���5��bV^{�m���5���:�>Ս�'"�س>�e\�ɘ]�1���)�mM�c�N�U D1g]�Ͽ���~�Ђ`��H�s2R���O'y�a\dh��m�,O���_�멒|���rct�S0���a�"X3h�xT9h��G@��GV�Ƣm���[W��f�P���d��O����F�.��.����K/K$�ٱ[��ރ��e]S������}�A�G
-�=��Kg[�lݺ�|�r<���������Iikj��~������in���L�z�Jvۛ=?1��� �+R�wF��|l����¤��΍xA�"ձ=\KTZ����(>��i;@w�t2I;uf@N� q�_��i���ad,��9 �CX)�s_/���ܜ��X�z��U}��9����RLF����im���*��*qۣ�o��V��ѷ�"�`�,.Lox����e5���Z6�m�W7��䆫k$ZEQ�#�28pUʺ`�T����2c]�i�)a� b���Y���-���'�K���އۈH� �� ���{cx.C�u�8ks0lbm��⬴Fız6LŖks0 �~-���AԪ��ҬL�)ll�}0�C�O!�a�@#��!�1bT�e+�ۺ�:�{�53J��5;ʘM�0 ܵ�<L�<85��ء�}$��i6�e��8��1�T� �_% Wȷ�$������er:��W�-]t���	I%��YM�9с�=��KWg��|����$R�)��vXڷ�"�}�������
�W�inE�5e�����#R����sIy���e�ޝ��ZU�������K���x�=_ ��h�����ȵ�=��_g0hkm6�>�|��r���
N<����������4��4���`���K������-R	H|q�j��7����@����Q_�ĺ,-���t"a{-�����ƈL����+�e�&��P��hД��=ú'�sxk�r�:��%1u||Q�x��膧��ȼ�^���gu})+�������>
�>s�2�
J�����O8������3�K��Z�v}X�����R_[%5�����rE����
�V�&1j6�?C&���&/���I�o|� 6xc�Y:�p� |���s%�@��`4*+�z��|��]����g�O���K����%���/��-�fy����W�(�:�k�{���ڱ^��u�����\�e����s�C�<�._�XG{���*�Q=�8�~F��v��&�fmϡ�W��/�*{v�fV��t�C�/P�D2~�uK�5�_Jz>,�(�|���laA������2j`|I����,ۆ��TTq}�..P$��X�e�j�%R������1���y5�%g^�[b3�N�lHH�$��0���4}|�S����&�ѐT�󟟖�W�r���
ccq�a���Eڐ�,�$6;A�[�PzfB�����6�%ٽ����PWݚ�9�ۆ�:G�NS�B�Ae�$�������
�S�<�Y9�ԍ�o����6�k`AlP�|pa�6�R `��66>)Ǔ�pt�%L�k�K�d�T�e�%�!�n��;lSHĝ�`�3��O��3~�F�J���r�?91��>5z�?9t��dX%��a�'�����rƎm=�BIY[���')�@�~UF9�?6��$i���^7|]�2�B�d�ԃrq~ZV�����S,���)�V��Jr���r��[j����C����<��㲶$ӹǾff&(��~�b����[�kʆ]��ݱ���a�	�f!�2U �k����f��q�m���m�`�є�6�X��Q�ƌE�8���헔�_ ����\"R���H �!��d��N:de��g�׌�NdWx~�i�F���r����FK*�I	����m� 6n**���ڢ�N1`��UAŤl��r��6&�,����'�Ï��w�ZcY.=�Я�)2�g��_����,���z�-���������y9{���;��8	}���*qil����+�8�H}����H��1��n�D�~0�gV�6���ND�$��5A���E��!�z���Ϟ{��Y�(D���q��������o@_��qr�g���/.��s�9�泍d�*�C�l�*�ҽ�����^x��X�9�=������x��VH�f
����.\�(�K��X+ �.���g�|��en�/��h]�\�!g�_%�R c�t�(�ϗ�E��*�B���/�Ո�v��nBL��?yZ���@��^q�J0�4�|�4�p�I��L�.Q��Ofj��iB�S�&�4�WG��a���%���j��.���s���Y���9�]�����S��2�WTs!A��r��jPhM�R��`��8(�*ȳ �N����y�������P��x��ΆV��j��~��aEƐב���^�?(͸�
<o≬����;��UAp>W���ڃʋ�/C�ϳ��͒-ŀ�%TlX}H��� ���(@/������>HЂkrx���'O��P\�ٲeP�-
��hb)B�q�ן���1ɂ鮬�'�*�O�me$���>o��,W��LϤ�%�zn�爓Da�&3����F*�B)����<�(�H�?�������60d��r6�	Ns�����f�T�	m'��@�l:�u�O���H���琚0_���mP�31J�
����0Z���1Q�9��PU5+�eR"4���eK{�\��R�e ���h9�V�+m���_���_����/�������(M�Q��q1c�g��2~�0�u���iy�A<[ �����<n"T�4�i����(fK�C@M5�hg%���4��K؇���fr��t^Hrm���������# m���M�MKl-.E�l�[v(z���C;H�k���1�p��X�d �O���%�q�y#���|�^0��|!�
~�K�B�4�U�����5C� Hk��Q1gƾ���3;���9Z����T�#c�����-0#�i�l4��IVMe�"�RR��A���<��<�� }�V����L�tP1i��ׂ�iѩ��	"�A�8���@n�y(wo٠����ZM�Ő�	^�����.�A��l"I��!�*8AFYʖXN��2腵�A��ڍQ�~֞��B_OӶ!�MB���x���YK�ȰT�P��-���L�������$	P�F�Z	׳�Η�4z�wG�>c\~C�:���n�:*�hؙ.8�$�op�������8��	-��:���u���+$ⱞps�PEu�@���A*7>+ͭ��Iba�Y�7�h0��5��Y������.��c*5Q�?�i@�9����RL������z�_�A��T�C?�z���1AN\���^7�S@A�`k�m|�������
�캮��7}fy��� h���ӠGR %=��'�I�����z31��11�b�MPC#�E'� ��h�vh����|UV�{���9Y����c���`uV�瞳��knni�l�F0>gS�q����`Dh$5:mr�L\���B;�5:Up����f���Xg���Sx6���\,�{�q�c�=� ��
�J!ں+�JUf����MG���)�*�&�m��� �&��E���իl+{�.0z�z6@��vf6��B�S���F�6@i�Jps�8���.~5HÔ)�!�R�1-��s�m�5�3�d�1cW5HX��:� ��d
�H���݅5{C�Uy�!��&.L�߈��r���(-[�[h��t���L^<��_�C��l��C�
�?� ��!MF�s2u�`��Kj˛�@N�:)#c+�D���� R����� !�i��y���9��a|~��g�Q��W��m�K��e/��8�$h���4�����PD���?����z���46x��-a��d3O,i�z�F3i��T�f\�ht��q4�A�2F�l�V������S��
I��t�h��$�p�N<)���&�s�o�E�f�e���х�hKX1p#�N�����X;T�Dv�2.|�Zx��Сԗa[b�+4 s�32;3Ev@S�Y	h,��|�aAY���y��3Q�ѯnz5��=e�83z�zԙ�kD��,[q���f�J#�;P!�d��:B����艢%��yC�"2;*j��K�1/U�<����4]4V]���lvj�zdeV����'��pBm5|���@�bQ�',Qw��W2|*�R�1��	�7��1)�s��J��21(��\�1I]`bF���b�*��f�`[q�@)9?ꭶ� S�	���,�E�m��U�1�vϚ� {M��$V6�� ��{_�z��m��B:ۓ��x*z!k�ؔg��f�~
���Tf�<ɻ��4F\,"H����3̹e��*&&�F�g���_� �����Jm�=�_!�E}���rB4�%(����$X�m� '�o�6�I�Dqdh���B�F}kC3=4pp@>7m����IƆ�i-b�����S�� �tI(,�g�2�#�_�����6c�I	��eRo:͈m$T�2�uD�	� CM[Z<	[�fRm:�@��s����!�<)��5rH���K$ �s&� �%3;�.��0!��� ϖk����*Z;�
�E�v�Z8z->Xo�c+5�� �\4����.
���}��c�MqmZ�m7q���U�0��jޓ�E��:�Q����S��h 6�i�nm���p�+FRMw�Q`�a�.mVjCV���d�iA�KM�PY�#�2Ft��O�
`�P}���&Z�sRf2FZ�@�ʎ��IzR�7H� X�咠];5���b%��Gؖ��j⦺0nޭQa�u��e��eӣ˧� @�j��'�L2Y�K�n���<�́���;;F��P���7�h��@���OW���(��6��i0��Z��O���v�j� %KfD�{ZF���{@"(H�����a\�O7���>���`�9��+6vJ�� �L:E~&�!dP����sdx@&'�Y���ϲ�*.�q�?b4�ؐ��bO0ة.��a"��)�B5XGO�l�Al�$��h!r�Q9򡄭E}OMV���}�����K�0s�jt��:�	ĄJ��f��ڜ)  @߿���(k07;1�Y 8N7ev8���5)+�t`�b�SV
e�S�Y˹�QQ/��(�X�,a ٦��җ���������07E�\!�*'�m:y���=���1?<��+@|�p�!�@&�Z��#H#7>����聒�|ԉ�O��O�.F=�&GҕE�g�Q�b��J���̂���13�ZՔ���'��>B+&�$��	ϻ��C�"v%�g��M/J���цS@<&ò�e�"������V����1��];1���#��B�P�q�:��0��^c����h��L!ǱY�<�p��mu����p�V!�� F����8�3�*9<7�!ZO�Pڪ\��\�����(�g��uKܘz�a���-S��#�J�|���"�}2d�ҹa�l���9{�~ޖL�u��]�o�#Ƌ�^H���Af�I6d������0��e��!c7�����w�UY�L0v(�f�����c�F51�j��	[S�������w3u�1t��`�r��A`�G�A�	e렳��F� ���`	��W@�<q:5�>�Ձ�I��A�?ÞV47
mT
���Zl	�-	@�)GN靶mu;���$+ �}���������Ta�1���W����	��U�/ƀ���^<wF�5�5���>���!_(v�S�_]hrʥ����3]�~�8z�v>��6L�U�4#ԽLԖ�SH/o[�INk�[�9u>I��m�t��Fw�V/�]5��`��g�1���r	^6�O?���h�����8���3 -^��@%ȧ)8$�1�ǂ���^��Z�K`���M$wc=�߇��oK��@?�����c[7K�x�v�>U��!p�c͆f����ߨ��p�����1\�qKq�t�E�^#깙Y����ܚ�Gk�Ed�I�����f��Uկ@�%K�N�_�y���s��IV��c+e���Uc+dd���i��Y�>�1i�/]�YFG�I�N@����>~B�NLJ�m����[����;yB���P�@��uV˦��2?7��f���\��*��kɌ{���[]��;$�N\�,&i�"(�L��W��Qc��|��Y�N�˝۷��Mdݚ1^��Ν{��wwI>,�Z ���r|�sL��N)]�Q�0���mW���8�@�w����Q��?�������Pt�B/���Wep=�P@�da��e�pé�l��S��Q$��~���YU�{�s�) l6r��Jwj��t�p,���w��srj�?ˀ͂	 �`�Md94ޘ(ǌ�C�(��1�CJ��4p|Q@��F��5��kո��9D5C̑��X/���%�{�1�ˀb3Ti�"i�5I�t�����-1���cl���6G.����)�������eK�32�<6& $0�G�[���eir�O�u�ZT�H[����3iw\�ᦗ�� �`��	��π��s6*���� N��U��|%l��� �{�ʆjol��(��q[���1Q\#�Cc��fs.HZ�����5��7??����ЕA����������%\���w��Q������(��0������H�J�<Jb
���3�M�k�%��r�{_���%��s^r��&�K��45!W#I-��S��oE���Z���
��Y�G��X�o	.t�@ۏ$B��v!�ڳ��b��0�$QM�F�%��JZ��"GJ�_	��Ş@������a�⪝�܄��?�x�?���	���W���T&�˱�ƀ��{�*2�:����ˁȣ~��~����v$I`��[Mk�t>�x����;R+�F�����'>`�qp	�M �ݢc�a�M�#G{�ă���_3�f%pV5�Q���@l������|����(ކI��j��㣏>�Ç���[�VZ�S�kM�E�D���>Ak	Xt���H|ݺr��[�7� r1TF8 ���9Ҟ����e����BV�R0��rO�-�o}�(�����S�m��r�8��J�ksajF��{?�_M�]w������Q���)f� u=t�ݲa�*��w�I
�����ɽ��)�i4�Z�Iٵ��|�{�*��[� �.��8ډ�%����_b�9#�n�&_x�~�@,L��zd�e�3X�p�i ���Y@�f<L<@�����J�\`�i'M�)Y���:�u�'vb�tU��ĥ�Ȧm�9�����s�*��Z�9�s�"O���\�E�ct��-�)8�D��h(�������Ԍ�,U#�B��$p `-h�D��o�"�)A�/RAn�v���$t�
�<N[%&a�j�g��Sh�8��M}X�F6R�;�؄�3��
8���v��K%���{)b���#вloi�;��#�87�E�L���H:�v�bdY���A�t�$+��
�O�Z�3d�(�[đ���ϽcfE+���I.2�Giܤ �o�颪�g�20ص���?�8&�82,˖K5th!��o��^���A�/�[)�P�MŦmR�՘���2�jZ�:y����թ�x�|pv�VL�Ջ�nE� �� �k��Ol=o��d�Gy�RJ�8��9I<+;{��@�n�̜:�� ��;�XlӍYW��L'�DG`��8V��a�;ZB�Mb� k��$��V,.{�R��,��l���}xփ e�=0�>��˲��Ke��*NͣBeݔe�����$�Aϵ�^'o����8wAv<�~6G�����ͷ�\�R(�����G�,ϊ�{.a�*[���?s�m׾�]"&|n=�b/�3&�:�k�ju�)���'�O�����8/���oL�K�g���Wn�~yQ���Z�s��R[�Wg���M���ܘ0��!Zv����;o��doo�f�Yٻk7�܌�6�pш��M���It3�Q�lFݚ�r�^1fO�8!gN�b�2��(�� 3� ���7�`L����`��0\�q�aLu�n�R�R#T:o��:���(�����M�u�O?��=�:���9]!==e^�!����~�?����7ʃ�����?��LM���e�X�U����~�uKz�Eu&c�%Y3�#7]s�<��N�p~N�_˙�����z�\s��r��7��,ZQ}�R���QSB�rUj��@WJ�|�RҬ��߼('O���e��+d���/?��>���\�c���:�
�g�MQ��`1l}I��SsB�M�IZ��l������4�m]�7`ePd� 1���j�jDN�:���a��jЧ��z���P#��SkC�V��a�j�[�`)��,;��N~���,�8�ny��X�����j�x��&��op�>kmy�<X������~�}�3�a�:�-�C+�Bl)E̒������4����'�K;�/	0"*�s,���W��m�Ծ������_�JÒ|�uB�2��t��ȍ��ي�t��������l%���F�I�:
7Ys�����H�Ct�G|E�3)S�k���Y���Z��a�ݢ�n����(�w�����j�y�Ue��]b�����"0jv�GP�@5��=k�6)��ci��,��cB�h5��<��γYk,N��Pp�ig�& ���vԒ���%L:$f�i,��V*�gl�,��Lk)Z����N��)Y���G�eF�I�d_[αB<���C�uB�|�8{o�h��M�}�� �А�e�~���~͚u��.���ݹ�k-*pg-�ͫ�j0@1�������v�||�����˲��[ȵE`�S0�6��Aص	�ޘ `���jM~�0tcA�* �Km{l��KJ�.����we)�h2��{�u I�Yg`��w���UT�(��F�0��� {�@ۣ�f�@ �YN�`���)7X��s3%,�4�sQe��6M��"� ���1����(:!ˤ��I��a�&��B�6�.���X�8��a2?7K�"F�8�8�3��aC���-ɀn�g��k��Ht8������{Y����,��{?�/�N��l�l
�g��ޡ��[*�y���`�^�?G %�!���{>+�֬�v�T�@�
8�\��+WIO1'}��y��s�d�P�";�xK^|�N���Ԍ�(׭��W]Ź{.���Z:�퓢�>ĹN�>)��9��f��I}aN�(]��걍r����O�|�)9�gu3!	���Ĕh�r!�_�R���i�*֣��Zw���q��tU�Xu �uDK��aܫ�Yj�X�#�r����5�a��p����x�2�HdgI���Ć��(��1���M�6f���Ȫ)��~:�@��=��-o�=N����gI�!b��߶}<�����t��K�<|�N����t�v7�I�>I��8p�E�V��=�kW�9_�#��&�\�W�F��� P[ׅ�1m��0���&f��'1H�����/�6N�.pm��2bD����t+t♎�"��X�ۃ�.�Au�eA0�7�v�pj��v��������TrN��C���;������c{0�<�Ό�k%/���I�;#�����X0�`���z�ЁA!	|I���k�����[��`?AL��F�W	�..��1���JWl��|0M�rn���i�0M�.!�e�c`iqU2�I�>���"8e&5%���6�l��Z���of��1b`�P�f���o��w�!_���������ı��jtDΫ�}䙩i@��D�ݬW�k�h��ᇲk�G2�b����C�k�z�����ʹ��-��<�0����f��A�Z�!�,"��2�;S��4P�Ev�boK�{�_h�002{�b8J���3�+�n�R��������;����g�,�������$3}�̐�FdEM���>��_�=�߰A�`t�h���	��9�0��3L|?�Y72�h�y�۝;?�2(*1ha|8�&5��p�m��覊�ܗ��hg k�H��գQ��������o�7)F""�4C��w'od�I��vFŨ�x�yzb��21~�2�Y�L�ªᬼ�ߕ�k+�[��D&E�$�l�dn�&��L��Y����'4 Ldhp��X�4p��G�U�!���̜z� ҥo�@�u��'����aX�f�\v�2;]�s�.���4E�2�*�
x۱����Џ�uxh��	pEk�a f��7�Onķ��`<�oE���I�B`���T X 8��wT5x�V�n�q���#P!�nj�O�����%I�D�1�l��됚/�L�g��M�������E\:<��Ա�� ȼ��
�0W鰞��е̹<[��u,�]�_���m=N?����|د�,���F^Mw�k��w ]Fi���(�V�ҝ�$ Z���RP*�tOU�2H� ���{�v
z�u���g��f�c�̨�UR��J�c���8R����zR�u��+��R�k � )YP8�� q<M������z (�����y��_b詊UR��Z��KB�b�D�SB��w��n���:�!�UJ��p�|���w�vo6%�v�D.x�k�vU��Z�Zy]!<��ĘXk3�$�k�;��� C�����X5 ��Iy����b�N\:oՇ"�*{�^,���~A��ve��B�J��X?m�*�ػuM��A�_��!��}U�����|��&G��H�>�T >�-	��R9�>%����܏~�q�r������=v�cپU�ې��,�|[ni�ђ�ĉ�~��.������ߴZ�p&ҭ������*^�b����W�b���kh�$�Χ.P�$��b2��<ω�s��1�87>N��J��CHb�٘='�s�%ٓ+�F~S,������ٳ��e��''gYb��Ԡ����n��Ug�0�L�N��������C����C�ʼ:b87������Q�f5H�7��ëT.t�0�G�j/Ď�+6_B`��}�����4V��JQ~�Q����������2���B{��`v��R� ���ؕ/�$���@�� fN?�~��N�����^u
X_48o8�vk�2>8OT@�8 �,ű1mR���I���y �:��n�]{�1��/�{��*S(�wX�AaU� s���D���V�5=��q����r��˱^v�-���N�$�v���ɸ|��#s�L࣌�Ybll�'�͓qX�F6s���RZ4����%�j��y�&(� b¸���$��A��@������'�G� �3Pj���ȶk�s��a�$r�襐@,c|$���˴�3�5�~�@g�z�	�6c*��s0�Y*��B!;��!4l8��SSU��1'0\)9q i?���>T�`*��씞����ڕ�&Ꙁ����0M�M��MG|Ȓ} ]�'Z��e	��=����~0��)q�� ���#�����)��9u���~VsT`�ρYtm�e����K�jύ'�<ꘃ���'�A��6���`U(pI-��)M�8��^Ck��]��G�kt�M�;7-��"!��	/����v.�k���C��
adD�݊�φo}��3&�Nh�VS����6 �:�	�v��tm�j�O|�7q��I��4�Uom#ǯ�I��A�4+F�I��ւ�rמ��c�g_p ]�6�x�
8_i��7�z�D���������������}{eQ��#�&���dʠj*&m����/k6��o}����3�8ہjy�1�6N�q��A����r���-Oq\'���rk���f��L���W`Ŵ�P�Ù��6&m kۑ��Xj����mD�7�ɤa&^����~[�J����� ��#�wg)W �v���!p�T��.�Q<���q�9YPi㽭�i5lS݇980�'�e�� =��R�3D� �s�j�v��KC�ŀ��M�H3v��l!GGT,��x�h�Xf�Z�!&"�Q��̬��� ��Ēl۶�Tۨ\�u���gOʉ���pi��2<<,�'�����vTB�DIFG���МN����ea~VV��}�4��e�'�` ��ZR]�UG=�m��8Ùa�C	y�
�U=���Z�Ѵ��ڢ� ���F��t�ONH%r�:�%r�gn�/���^���>'/��*7?���*`�;F�l�(����A@�(�B�N�U�rO�*߇�>�n��g��=�����Of-r�����"�
��ol�q����@Af���@�Qo$x���
E�/y#;��k�N�ݓUh������P7���f�:.���oj�B=&��q.�X_>��[yGU
�Fur�f`j­���s6q���{Z5�[�T�������z�ih<9��Ъ��`��A��+9�s� !����$�V!CP�$}�2�A�}X -�9�7�s0q�g�Ā%z={�-g���a'�̡�Ծ�;66L���)� ��IL��I�����\7t��p9��Ǡ�ڰ5�ʛ��\�նذ���!��[G`m.v�y`��L��\[S,s*�ۄ�L�k�&��%�}l�V�F`���RR:`' &.p�� /�-��e��Ct��M0�Nح8�rdSu�<3l$K<�ƃ�瑺�ZC6t�`sq�����^{����c\W8G�	�Եv�t��*�I�q}^-��MŃR�6�뮢m�h�5w��J>��"�~���)����U����{y�Oɱ#GY5F�߹0;Gvj�v������Qy����vIC��%��L�Z�7t��H�b?y����\�6���%f��5N�&��`]�����k�9����%��3v�q}Q�׋�&c�$`I���A"��z���6Gױ�Y9;~Q3�"A�5���˼���>3��-4�j"�J`��R�nB��o؁���ߝ���V��H�2�����K~d6��^����v�� H��'��3	�^����3��\/0`�v�B0��Z��5j���檫6˟����'����Ց-�/�/�zJv��O�wh���F1���&�^=&V}�,�����Z�_�J�iP�&�� ʷ��r������q�ܴ�F�x���744L�Gpu�@�I�T�\ew�v*R(u���]�)����m�'cJC׺�'���ؔm7])>r���X~�'���_d�DKa�@=�01�5�j�}��)�aj�4C �S�)5^K��1��g����r��U6���n$7a�-�)6�i졑+{�~A�t��I�A�6�b`N_���B����Z�\�����@EZ9�%�{��}f�<�m�c�{n�@FTq#��rA�b��]HМ�ZPݠjb���(�֔��*�2k*F��@�ؠҵ�

p��RA��a�<��a&��yp��,�C���Ƞ"��	���\{��x�׃�����	UD<���)9^[��7�� � .��6�)r�֛�z-1f70n����z��IW�@�I�ʬ&��ܠZH�����P!��ƺ�uO���g۩�u(��Yq�2��n2����}W`N����TX�" Vo��B��8d�F�6EH�@ώ�"H��qmbih`��5��@��_��;R>c,��̔���V� cp������$:��9�S���Jnw���}�K8��8�)�Lg���8U$\�2k� v<F,�a�TIqm�-�V��p�� �6�3A�xn�ݭ�5��sQ�gyRmM�6c����|�Iǋ/�!�S��?��?�_���;	5K9��8�j�IA8ypv}�[ߖW^{��A�ܯ~oBz������9k��3�Lp�c��!��W���� G+�0jr����Ib�*�1�Z��"c�0�3ŞG��E���X}���������i�OFE�}�AІ�
� �i�qQ2+m�	�7<K���K���7~fP9έ�f�Y�Mn�Ao9-`�d��j�9���4(�ˀ���ܩS�$	��X�B���=a�r+@��P��ʪ��\��ae@��Y�x?z�`Kd������r�m2�j��J%s��>uBΞ9e-��@����r��Y,̯�w��1-�e˕r�9��qy�ý@�.�|��|���?��?�'��]Vs��+_f���_���Y���:(���!�R��k֎II��.���C ������>�����d�?#��{�|�K_�Z�_�#�������i͘��-6\۪��������>�F�!f�@���:��x�nI4pc�"��2�='���J&��K\vHǎ�	}� �
�8u�C�q!����?���k:�+���-����' �k'm�R���A���c\-T�ă1��!{��f�ВB�x���	@YR��Uf��̄br�dA�nՠ�5�a_Y$�H_��$:=3�ԫ3\�lP`f��c�Jڎ���J����t�˦�\69q͎��6[\z(W������#�u�ԙ��`<G��S��]�u�@�A.R`'a_�p~:�=�L�*��B�-�05�4g	�Xrb��ѸcD#T[q�R����?�ʄ�I13mV��Mft�7�t�|��b҇�ĵ��rA
*#h�EV=N��Wa �jtd~v��b NL�έv���~��$�q�5��ұ�.@Ap�q�@d�pN��/�~`S=�+?�
�f<��+X��9zxgwf�����f��$�2�^U�A�#�� �]�E�0%n�(u%ORHVV�/4y��X�E	�a|?3I9�M@,���n˟Ľa�����TR�:�����Ͷ�]����!=z.ʃ#r��9�O���*�߰�g��H*����z(nC�h||\�/^���1�u'C�+9�v�W�;%�Ă�k��?��pq�S����^'r'�� ���N�,���jS.�:��X�+H������E�r�|�xa���%�&3�!�����[O�[4��f
���!Q�Ԗ1dC����[V�B5�Mr��Vn����H��H��P�1R�u���}^�P��`Q05-���� k4C��K���Gmb���J�ņ@��������p �ѫF�����Ǐ��Ȁ�x���z�z�Tf��R��e�txd��^[妆�p4�wh���KA���'��O~�˔���+�~�1��}w�řEy��'%T���3/JK�C�-���?0����o}�	y��7��s�U9{aA~��/I^����l�����d��XZ(��,�T_��&�ɭ�ׇ\���U���ǈ[y������\s�V�N�<����_6���~'J���\�0.�^G�� �+��S��z#���d,��8��L�	�(N����M�dr]t?��]� /TQXM��t:�@��Z1�j��,!�}��K舐��j0.�:b�3�]�[�,�$t3C��јā\����ǻ,�A��(`&	.��~	*y/)��22>S%سOT��{Ї� ��֭�A����c�4����u�e�p/����<'�(NdxhL*=%b���B�R,��Az5��8��d&:-w�mj�X���`���r|7����Qz�F��T����!F���F�65���*�<�֖Y"��L�[�#J��0��f]��ޠ��vRªXL|U�A�z��f���uq
�h�ږ��%��Sb�Al��ʆIŎ��6��Ṁ'
l��C�#:�*\p�<�ْTu�l�������������>�N�4p�a�t؍�7r�qi��8���l���Wb3<,{Xu"p�&�Z�;V/&��*�]K�`G'>�wg����>�WE?MB��t�8�D�s��T�擁:c��ā��l��WX��2���#�x�Ħ��t+~��Rx��M�r=ȳ���2�6v���/�z^}{�K �)ms����8�}��7@�1E�/WȒ��\�c0�W�ߊ�� ���#�m�9QX
ց�K ���u mK�M#~4L�|+�qV�ho,�$��*�1�R��g�<�Cp]���IҚ�<��L>]���s[iR֍�{˜L	\i	#*)e�;�1*�B0�I�d��@�FU3���S)�MqА�q���艇��~;veǔr����aɩA%a�`�,+ �ʑ^�E���cTDI�DD�Au����6����zj`Lp�]�:uJv��!_��#G>66*�/��^yU3��̨C�j���������l�Y/��v��)~��jr%�5�P�����<�k�
_�-[��{�Iu�O��W_{�Y�wl������Ev��h���S�v��o��_~P��c��c��8������4�^�J�:ƌfLø(�s����4ۮKA��m[���@E��D��|�|����`'�)]��_~Y���3\ë��J}��v���:cu���c���tkr�=w��;����?�{���ٜ3�n���ma6�&}�&vH�A�,����ԕ��3���'p���o,I;����H��1,�B4�4��CƤ�}�qI�8���=��ܨ(�_`:P�m�2�,�X��⢬Y5&_���r�UW��aj�"�+�H�̳��ZlfY�U(��G�[n�nmж����:-/�1���s�f�~�^�c�|Iv��#y��7�V�r�e�>$+V��% �0�_��d��t�ub<�e�|�@��y���ß{@ʅ�>ء�z+��U7������sr��	y��_i�ԡ��������x�~��ɫo�-u�P�!9����Z-�n�n�
�
��9�{�%���T�zeU���ɪME��A�ܘB�r�Buh-�X%��ǁ�Q�%`8G;E�zuj ��٪��9��S����ROY�����l���O�����|���B�K���!y�?�~Y�8$:�1��=J� @�h]Z� �*
�z�13�Ke¥]��4��e*��!@���ܛzg�7]u���R+��?=dՖ�"I���F�}S;�J�ϱ�D�|��NS��-R�G�s|u(�=��oSG�F�n�d{�����Ж)���9��Úq}�E~�(���Ґ�bת�|AT�0�����OFe�1F�(��טa�t��
r��
�ޱ��F�ŵ��{Z �jT�v+Z�Ӻ�mJ<�a��"4����Y@cd�1'@����קK�0\N���
�,�c�{���V�[d_` D4�L���DkA �Z���"DڨА� �Z�/��;6c�殒�����F��^_��Z�B⻯��:�0;o�����52���4�h�yP��6L�f�����]v�e�6S7���g�>wV��t#?����ߕ��#ǎ�2t��q���ϑ�����ǚ�z�>~JΜ������s32[ÔLF�:)S��Y�j��-�2WMet�F9{~Z����/G����I�����`#�S�����/�M������l�}��Iٻw/[G�r���G�c�h�!���}{v�s����F?��S�f�ãbta�9x@f4 ����o���>{e߇��!���͗ʎ{��ً�ȁG䋏<"�6�L��V�E�C�Z�v ��)v���h��{҉���� �v�+rA���Q��K7~	�~�W��Qx�(/#�$Dd��X�-�[�5OW����Q�'˩:5�F�,��@�k��6�]�l�UcE������?*�v���w�@MT��W��m7ߤ���c�8pF�>$��s���#h���\�0'ϟ;%��1�65yA���ի�5iX#O��9���`�rl�]v�,�hh�X�]�/��[)���Ǥ����=���;zftO���t?��S�9��Q��	Z��%�l`U�b��}ӹ�ڷ�PIja�M�>Ơav�󊱙�8�<Rj����"��v��쩧���IV}���
S+t�,+9V��Գ`3qkpD�RŪ=��C� cҎM�U���FR�N"�%�`��He� ֭�>�ѼhPj��g�#ŉc�EKݍNs�UWP�-p�?V��9�C
�hK�����e��2���0*��V#��0���g����7:��r�&W��SqH�3��80'I��0,���!��vm* �p92�XN��A��J��t�|vRW-��} �Ĺ�=�6����T(q�gv�ɂ��hG�ڏ �r�p_1��ȼ&��Ujp�@�(A������`��Œ&�J�i�a�;ւ	�@n)ǁ�I���]_Ib�)g��I�%�fo���h�M�l$&���p@�{Ej}X��02�����[	TP�/k��7���\��ۄ096�k��Z\X�04RzJr�$�>���K≠pP���8I0 �������sg��B  �
E���a@h���Ǉ̈́h�7���	���~Aehm�<y�n�H�m�$�O�"�	9�bZ��z�ȅi��r�{���򀣄`�Q��¬h|rA~���АLk�-LFe4S����!)�ɻ��骠�{����Pv|X9��B]7{>�*��^�Sϼ���S���T���d�-��-���K�3TGF��/Ԛ�LOO�1-ɶm�rM��[�p`�H��|��{2�V9)���:�Af��#�uC"�)�� H^��_���H�x�;r��)ٲe��r�-��$�C�:;(5�hW�����8r6*��@�"��C�31q�&ơBl�S��ُ+�@����E:`U+Urj(�8���CO�!�"j��^oؒ�qu�p3� ����L��BJ򎍁G˰6}�1���o�%��~��m���깩�lX�J�֠��S�6��C��ڭr���da�Fwa�&.^���sR낪I����Gr��9y��7�푉��䃝���5��3�m�׽g��273�ڰ9jpy0]9�Ǣ�W.����Ӳ�>Y|�~i-�\�����o�c�RW������?�c�x�f26C8q>��g�"&"��uu6���H��ԡ��M�G�R��e�سLnbk�R�����*�������8,O��Q��ފMY����-�?�����B�Au<`���&ZhL�;��!������[���\�cUvX�qM&0U�r�׳v�*b��f���g�Q��%:_{���|0���@�1��Po���rAM����с��
�{�[�cd�k=Z�΍��3�pY��	M�.q`Vb�2���a/���2x��q�$�r��1�Θ,���G �&c��:.T�}{I(&;���[5��t�+�aL�Ə��m$��l���"�K@4������@U8�cD�;2��p4��	�)�*~j��6���&|�����KT0�m	m ��{��Ó0 tk�j2���]�݉#yb&r���ܱ3��#&��Ւ�[1�M�H=�f|��*�Ĩ�`�����S���K�%N��Ư�J���R>SزysP.j�Y!�L�:�i���׫��0[%�B������C2�r�S>Ч@�JN��U\� ��c�r��q���G�a��c�j�x̓T�qu����9�n�@���:|
�v�P������!Y�F���T���Le}gu��G	;��ɗF��aPM5�Xɍ:�0��̜~f�,�p$�!�B�lTӓS�ݖѿ��n����^_�oX�	���^����h\�RE*�,�zf�fXB�@	�8M=H��\Z2W5���)��6da��� ���uy��4vPŝc�bfv�����ʑU�hv4\��������7�"����ܬ��]6y������,e�b��A�_��O1Ǚ�	����aP*�ïi�Y)���#M/�� ˒{D#���e�!��6��a�7��{g��>�#�aw�τ�Rfz'�kȚX&f����ǈ�q����W8�:
w���K� b��@{%qΗ�f8H�
�:�=�׀�j����Ƽ����������}�X�Vn�i��<r��P��C�]��֑���ET�R\3*L��Z�"� �JQ
��-��qH�7��01��� o�^�5��s�I���^�Q�/�v�n��yh��By�?��l�_dຨ6c��(G�A�_.[bG���ң�X_�����~��u�)�鎼:��z�����1V��«�{��͛�O���5���3z���e��C�@Ŧ��Y�1=61~^M���n\�^��?���L�h�x~���d5q��l~�.�^��^Y?ܣI��]�~����j��{�8���f�*9��G�;��P�뙓��чѫ���?22(×n`��V���L7ڥ�.Q[�˽z�����i�W�����T��kR�%Z|�)�L�"�Blk�� a!��s�u�0��q���G�p$�u�
$6rB�`�P�vZVm(��A<�Y,I(:��N�F��b�{��2��0�I��S�g[��V��p�ϑ;�x3l$����	.���_�q�Ё�Ѣ�@ڐe�g>���
O'�
H@��}n�P0�P�����sX����'V*��o�!j��1�^T;�&!���$�B������ւ����8��2"H���f [�dM�7&i�Ԃp�_T`���@�vuF}�%�9]�B.�ĵ��5�3���?���������8+ri�B���Wc^�h�s5ۆ �b�U�W�G�0� ��n*�fm��:�f�� c�
	m�?pV՚����g���hP�K�V�/���@Py�����cf��	^J �֬t�I�}����9uvRX�L�,�$*#(c抌�Q�����lQ  ��IDATibB�A��٣�b.�A�&��}L{ �%��0�`���MC�]�cy�2 �ܮrmH�0����,J%�+� �r��[ $k�S�����/hP�(ɞR `��T�r$D�����=k+�f�C�2����\���������[5��>a�!ȵ��N�ձL�Z2tod�}b��je����-��4�F
e}��F9SW=�e��J�>v�L'v:n���{uG	�hj}c�S#��t�>���F 藪���ŝ�*��k 6J�=�w�*0�'��f�T�nGrɦr������ңN���n���!y��W�$/B��0q<pLy�-ӨuȤ�箇�Z6�{�F��[���g+��l���7��@��g���:LL�poj��\�bذg�(q떫嶻>#���r��yy�Oʙ3���3���B}�qT�����Z��嚭��+���kײ���{�ʳ�>��������#���[�˚�kdT��Լ����%�n�" @����	��>��|@n�e�|�[�$�7l�;A�*��3|�]w�� ��������K�a�:����R�k͚5�$M�L��W�ʾ}Q�c��<�c�l�|�U�p?��UkV3){�7�?�>���o�?��?�ϑ9?��s���o���Q勏|��ۇV&0/�������A����'�OV���<�v��'���w�n KO��2�����K�%Eb��a�\u۫�0$V��B��\�m����J7?���&"�ͥ�Zʊ8� *,�~T#pC��fsYN�%���-�Ю� �/#h4\�IU��ψ�I�����I�//=5 �.Q�$���-��$6��TG�%1vs;ˮ���ua31C�vt�(��� ��dm�����Y$��r��5J��n`$�D
P<�4�ܰz-������M�՘:>���W�<t9��c��BUZoB/�q�L�Ks�dF*�5�����o�ǫ�������RK2�\C7���<{Ľ�A��:�iu�gf�4�h�!�q���
c04:d�6�"�i����aHZ|h�s�Z���+����!X��j{D�hy �_I^�-%Z�Q�PdO��`�N�E�ٷ�Q:vJ&ff9��L2W��<�?:seS�^C#���M���ؐrbb�.�?R�(+^�g$bDhjHt��13��t�]ڨ-�������Pa'��`�0Ʈ�= �u�()i�7���	�����c�J�pV�/�85���J��q5PBK���� ��	-��Fu����V��s&EPz�0��Aݔ쓘�!�T�S����60�Մ%��鸱IG���J�\�8����y��w�nv(�?��-���k8���z��7`���69�##�0uڔ-��S@����Z�:~�B��>yB���i-4eL3�{�$�K/7u�3g�8"Ec��/z�E��t��yB1�{��
�b��ٚ�w�8)�8�4虊kܯm̳���b	i9��k������=��῁�z��˯�J~��F��~W��{�3�:q$�}X�~�߇~D�9"/���r�,��@�|�k���|����?N�~�G���|��|�%lٜ<yܨ �m���hI�<s���pR�6�g����
����
'�֯]#�׭����������(?���p������ş�������<�A�YN��i�z!�V��sr��8?sX��n�U�����޽[>x�}������6I_$�&gҦ��������ߓO�X��^�~�V�������?�G{X��l�<����Ç�s��w�}�|�{�ѳX�>����Gr2�P�(�����S�������;%�����Ʈ��N�+1��8ε��f�VdP� ���L}�N��O���}�nCOV�ώx�˯շr}5d˨E��
*Z7�Ǡ�ˠ��'q���D%��|�3�.�b2g	�����"�5��>6; ��;�mۮcR�a�
ڥ�O0@���@��D ���U�y!��ˋ��	<�Aչ�����rH����<$��#������HR{{�����s�>�ǜ��bF ���ڵK��:yx��i�6a�{���vZ�Za^fNf5��DC~cn�TkVebzBf��h�X���Ypu��7������43 �Y�J��mv�������u�jp�u�7Y���HJ��� ���D;p��r-�[ufV��<7�]t#/�q����-x��f�6�̨у"�F���$3�e��e"�>��R;s\01�#7ph��aցB��}� �&(�UeN�pkCY��2S��J����3G��3� �]��0��D�bG�����reO���@-����)j�[,��i>*�wi��d�eW�#�<"�Μ�߼�3�0�ʙ��1㡇%� .c�_��y>j�`�;6쌕�Ǯ���%��qk�v�v���%��'f���a%��������p�����ggK�ҽ��I�F��oYZ��9=G ��ٽW>>pP�ٶ�Aȥ�o�~�Bp|����\ԽH|U�X:!C"?XP�-�����&E9*�gF�,�_~�f&�&lEy�80L���� ��>^�6Xڧ��� �u�ؚ׭[#[��Z�~�19FFV�3Mژ1Q����5�V���Y�z��t�R)r���:������r͕WȦu�Y�@v�Ȱ�߿_^z�y�����(#=���+/��>T�~)�mT_|�9p� 5}��NMk�;"��99w�%?��ly����d�ʶ������՗^�(��ӧd��ur���e߾}����ɬ��j5��y�yg���7�wt^��A��]�����t��8�d�	��h-�~�-�2r�����[�3�f�ub�֑To���u�*�}��|���$�����*;3~���|�W���1�/F!N7ޏgV�.)�P��IؒgK>y~��!S���X�i��MF`�)&̅K��E�p^�­��F��g����.M@��H蕟���8ʜ�*�]�q�����
?#�<�0�n|^^��8�4��P��&�lH`e��:��1qM�v8�0���ݱ
���U�_N����繟ZB������꽣m�rŰ���:���QFSn�"C[�K7�=w�J|�{�푃G��F&�
{U��&}��̹6:5��|����n�Q�z����N���ON�����a���$��<x��W��0<��Y�n�:�L����������!��usf�o�B`X�<D�4sDi?G�ߌ�Se�$M�5�t���d��i�[Aa��,��,�����l�f�y��i����+��P�� ;~JN��H�IV�Y|�Gt��1�w '5��+5eZ=���39lK�ʃ���
 �$����%2��S)7>^��q ��w�(��s	�c2�$ZG���UI��< ��	�J��)��߉��Z&�HdcM�eu,�Q�m�w�sA^G��C�Nɵ�^'�g�NeN֪ӹJ��@�fȟ�O��c��O��� @�P^�ӱ��]V�g����c��b��&9Z�@�@#�c}��
�hu���@!]F��N/M����r`�Ќ�X��UW�$�z_�3�[�^L'�aL�![ 8�=Ţ,�,�Ta�|��	/�r�U8�=r�����
N���]:�zS�F��r�K
����pL��0(ǎ�`�������E(-7xϠ4G�353/�Jy�PIL�':@�ǹ�,�,������ӑP0`נ	|3�N�9�[9�~��;���a#�r���;�^r�lڰ�c�c�+X1����7o� 9��'�1� a�_\���?f���'�kDu�����|_�{~������~F���L�}�gdT�j��βJ�V����, ^��Me�{;��`�<���Ej��`Ȕ��~����O��B�����*ק�I��! �C; ?Gˋ8�#o��&�֘ *eӦ�?���I���O��?����� ��g�B34N�n���r�>�����^Y��*���*M?��8���	r��������FvX08�0uAbSU�U�0��`Oǂ�D�փ�M
Y[�ˀ�'��3��
Jl��@
�<�=�e[I�)��y�qeG|�m����&�K;�"Oz'��Ӷ�]yN��Έ(�A2|؛��"g4i�:��u�)�����K6I��@��ԗ�6�03/2P�.,��<~�|�?����+o�#�k >��1̸�h�I���'Ӫ�Q@�53G�@߃3�X�	=��D���_=*W\y���o?e�
Pz�A+̆�.j��<8�]���1Y�\ӽ�� *�� F�,k�#Ռ:�I33+MnT0�4-jf�����Mf��n��=������.6� UEИ�͆�\���jSj�����)[��\��ƹ����2������i�Ku�-j.8.��ɴ�0l�tR��	�9ue�c|!� ��0Z��%GcY������M"�CB�O�$4 ^)t��T]u�,`�͒c"�a��\ll0f��ބXY�y�N ����qǜ��ŭ;�(���߀Do�Hj�M$���9�������|Y�]{=��V�.��������	z޴q�L�����\��jy�WY��t������ـϣ>_U'q������:��c7t��{a����o�~&Ŀ�s�Y�#�Ǡ�',in,��sj�jI��<|�����f�"�vf��*�-�N�l��w��a9p谬&F#���Kk*O��)9}�<��!�Ģ ���S��ڱ��=s^��X!8z�����g�ĩ��ӯ��|��ǩc�}Y�`B��� 0ŵP�<5�n�	��	�U��,�z5ڠ�$i��{�5}�w�}7֍6�)�'�ӳ6���[1�� 	�Ř�CP����]Wl������z�M�)J�y�5�̘&�^7:Z:?��S��#���.NN�-�r8�K���hK�7���/08@ �*8��w�>�{A+�m;,��2��u�B�L���d�e�Lm6�ѹ�y����Gy X�;�v��uJ�V���w�Zp �L�'L��s_}�5yp���Q���>��ᕣ�CX&P��@n��/֞ό+����(r��eUE۞���|���I�k�F�"򨠊�ɞ�U:q�E�ώ	&'�*�c��d
\����qf�B���]�t=�*<�*-.�"D'c
�"�HU�� ��jB���A�H
Rz*�[�:vUq�L�U`�`V��`p��.�} M+ufcL��tm�l�:ٴn5�BA6�c5�Y�V�jxH��NK/�f 9������j$��yCռG���P�����K���O��{OW]�4P9y��=}Jm̂�MOH6�L��iR��Ӫ���=&A&D��� Z
�yu�hKH��"�ACC7�^I�u�`�H���Ĩ��h�`r(��Ɖ5#(geaz\����
 ��ll�>{˕�!ӎMo��]��R�ڍ��뮓w�zU^{�k�X%[�����y~��� lK����ǭ��_�x���1Sc�"mR%θ�V�4�)}��+4�D��ܧ��h�V�g8����0o3���靐#�3"R���++�!�������Y�MF��\�
bG�ݘ���R/Ց�{�����!��?}[֪a��IG����#컮Y�Z���_��)�r��Qf��ͳ��kG���� �s����j Z�Hň��p
�%a�zr�'p���*!����r�:�i�ǉ��Y`(�Z�|bd9I}D�3N�S,]�}o7X�%��$�AO"��·��I��9P� 0Յ��yij�	��3����w�=}��~��gw��ٻ�c�I�CA%1¤�dx�,��'&��VC�h-0x�SG��@��1���aOFO�~�R��sf8��(��Mt\	x.�����}pLw�)���es����`:x�0 +�����t�p�p����J[�Ⱦ���/���a�&�b���\��sĨh�@���NLMr���q�-����Nd�h5B�]آH� �U�\/T�P颮 ��E�ٚ���V���9JRH@��E։CC����b�����#�T0o�:��&���1?ˠj�ƍ<����u���P�z��i��>�Ҁ-���s��ܵG�v�YKO�M�� '�X�������-l�+��`I����>�r��em?��9��3�O�%N!~�	%q���������cR�W��K0֓ �js�Gq��tϡk�{P<e��><�y+-�BQ2`�����U�e���pmݐMl1�� -u�T6B������6����qY�z�l�q����!:�\�IF��:7!��u��9� o���-IF?����d��zt_65���N�9�?N:͚�5HY9<�>�L������f���y)�~��{ � E��8d�y������]�t*��v�i��� ̗����'�R^6��,�������5���l����D9/f+����H�H����h�Ûmid��`���[Z�Rr�j�`�N��h�ѐ,�B'Q �uL>����\Ŀ�d��A��w�a	r5�t���+�D�����c���y5M�X�V�!�5�E���'����4�b�2�B�>���@V�J����'��h6)˓z�%#σ�A e�US
������l�ի�8a� '�vK��
��z6k������c�:��'OpmѦ*d��c�}9L�dLۂj�-9�>{�dc��]+Wn�Dn��jN44pɒ`)���ݷ����!���.�jP:<���װPgi���#����p�J$QZ8�?�nP�U|�Ě/��qYXjﵤ�[D�����t��삓.�856V��x���ʂ��[G��:�'Nܰ�7!�8�/��r�G�ABGZ��:�ɩ�p�^���;ex�G𼼷k�?}�gg^�͜:�{��,Ԛ$L�m����4f'����a�6���cI�R�7� Ζ{)I��vHFrd|n���,2P���-,<2Я��Ƞ����{d|zZ�s�,7ݼ]6_q�|���0U�b���,`�0�pV��M�o���Z] �N�Op��){xVvqb��/��s�	�S������-��~ܰ��䴞�6a��^u���/�L��	�0H|p���? W\~�P-@+��V�� `��;~q����څ	!��`�6�P��>/ꔩ��b%��3-h8q�lݺ�6ktlL��.N�@QA^&��ҧ�SO�J<(�<���[�b��&�u���s�]���������U��sU��s��f�?9�ij��s��)u}b���p`�3��821�8�UeB�JďNlB�������	�n��+�Tv|��[r�Sf��T��{�.�;l���BIr���6��b2
��3@�h���M9�<�6�(���.4ψ+I��j`>�����WΫb�a#��=e&w �?9�I��5@�9#6�5	MG����5[���>��8=���g��DU~r|����C�zl�t�Miocj[��<;�9���Z%c+W�a�������?]��(���TC�v�K�ʶ�����u�>�(��=�Hz�s������Dv����A���OA܄��:��|�\��2��������W4����������1�U쩘SIQ�(P`-%����'O��={hr�:�-�8qꜼ��r��,3- ��>�����-N�74@���%{��X 8e��6fh�^T]8n��"~$�� Qd %(q泔7n�D�|��jvLap�J�G�y���0��]"b�g�~�!�{XuX�j�l�M�ߝ:�S$̂Qv��hƯ����u+Vh$�O���cG��4��(T����K>�;��6Gq�0��v)�A��T��W�dF5��TB��rq�DQ�ZLp����75T�X֍������/��
��{��bX��**�Y�@�W0`���J\y�W`�<��1�=O9���N��߂-ఀ��.�Z;���M
$T�]�z��CC�2��s�VD�'�Q�'O���ݛ?�u�gb�9��[��h4� �;�E�$��(Q���L��{Tv<��8N�J���TR�_2v�L�v�%Y��Q$E�� )�7�w߾�z���<�wn�g�'ZU�,�^�=�;�����<o�}N�g������IH��l �(y��B��#��C(Љ��QlL���d1�32�q��#h�>���t�L�h�X�#7�ؤ��.�C����F�:�w�T���aw�/W>�&�)y����}V67�y/p��BI����-����s�|f[&�[�O>��s�w?{M&�&��y���r��uY���*MϿ����jr��+�~���uppv��
�919MR7T쀑Z8�D,˦(���9��;�weW����,��h�@�Sq+4^��*�90��{N���k@}1��@P�T���C�I/T�0مd#��5��g�e}S���ѣd0B�����W^�����+\����Pb�`��A������ٳ�'B��޾�Bۈ�<N�����h�:���q�N����pC�	_&�u@jo��f���I��~zI�{m!~��^q�wv�&�h������i�Ĳ�1�6��"k[�+����Z��-A+X�n�%�Q_
8�Z .�msz2���g�+����M�n~d�L$�j�L���+����aטׁ1��6��F��II�(�� qʥ���d��AJ}oK����:M�oS����=ynfR�]�<%+?yYvw�	?�Z���`�Qe�(�ק��PH��o���G+Uҵ�h�%�ң�<�k�	�I��D������OL���nr)P]�kX��)��x�@ѻ>��QPq�����VN� �S7|6�҃VdrW�H��u7{"7VV��qseU��� ��R6᠟��I����@f$~�)�:����r���r���M�o��r����oB��J)���҃���@�yw@"����I*&rP�`�$Ѯ�@����FϺ��$$E؄p2Mu,F�,xH�e(�,��I=�@��bS�D��0���ZudJ�xS 2e�*�~�YB�h{<��� ~��m�~$���ɓ�<"s� nt|�f�m@"i��<HC�(���739����]�!o��v[&��ƣ3�ɩ2+,m�=7`��c*�˨:$��Hַ��J�ݖ�ů}M�/��+hIe�1#̎�,e|o�7��L�������~'�,k�N����C�r4���ȺH���H�q�p��I�3����]�*q����r���&�&��_f�cyy�:�4k�>x��yࡇ��X�X�����Ȉ��S����g	�����9B���2���#��ڤ�`$(����en��#�#ހ'�f,0��/ex��"&����8qB��
A���OȒ�̢��^xOj��=�(�w�C�ߖ���{����srJ����}�=_��W�a��j�}��˯�"s��>�������s�����/#�*~�0����,���/�[����~��~#�A�qqq��@��k�Z�����^`AV��h�" 	�~�C�8�D�&tc�G��ʄK�t�p�|���9uVx���`	���k��*�>zF������YA^[ې��k���b�����x����m9w�]� �1�����% �X�3J�Q4�K�|j�&!@�ql��q5cLU��� 5��1}k9<A�#V��J��.RrO(����������OÕ��,��E0!Y��)gc�_)pb�P+��	\'�(��8�/�A�x�Pm�`� g k�2��	C55QS%�{]��j2��w�"�����*��Ag�@�\̒M����H�:ͦ�LO�ґ�d������{Q0������/&>I��nq���~��q���uW��^}�R���v��!�ӠG�̤.�(�h4��q-h?��N"�q� ^��q�ia�Ӿ�B��d$�r��j���02�QPc/�><��k�W�g�8��8K�Љ�ث�r�i&p��G�z�;����e�d�d��v���ߘ� �C:N��s�D_GN�J���[o�-Ͻ#E}���_�+y�Sgz��Zc���3\�@7��������QQ֋ݨ����N�z���S<��ز	0���[��>�[U	TL�U��7����R���顪V�������Oq���f{���Eڗr)ER�>2�����"3:|66}Dv����+���H���){�m����:zG�3v�\
>��:�`�+�BZ�Vnȭk����Y��TI6's���� �a-�j� c�I�H�´��޹*)}�
J�Q�T��g、��ͮ��7T��C�!�S�+{x�Fh6�J��rJ���눠r���p�h �񷄤7��XU�ժK��]KIdܘ�8�xK��ʺ�,"F����QuL��t`z䕟��1\�p� �ĸ2��`lEka���������S'������AŐL�SU�#�`Fp� C�wA0������}��	�5�Rȉ�|�̫���e�ݑ	�/0����3N�>-G�.I��#�ŋ�Ҡ�k]Y����U���k�l��^�#>�0���~���˅�����*���_��>{��~�4�ՠs���[o�A�����3�<�������9f�௸~���u#�C�����`��� ��;ߖMv����[S���@.��K��ٵ��ׇ@��?�!��w��eu:�n\���3a��4#&�S�㇗/irw��ܨ� �X_�����Nϙ3g�"���{��os�Ɩh�i��������j+o��g�|]����7���)ND����B�A/i�~���״k�2pSr�= ��Oh�43N4�B;���)���}QM�M��������C$��AR;�F�i6�ɢ(v��F���S����+��"�U����~`QEZ�{�V�ըIQ�8p#T�f�.�%ة�^�g"pM�{e4�4��j��6 7T�X��!YTv�74(YdSf�X��llm��
&0W�|֤T�y=G��Ee.(M>���P�C��3�8L`�����6���׽��HmcC�@�qh��P9��`��k{}"�JN���tLI��#7Q��Y��z{!�&��?�oNJ��؈��W~cd직��x �@���������dKU	�mF��������A�,z�i8�l�=�>��f��y�
�x�xD��{<Hц�=�/�NQD��ћ���
��㦝 Ud�Qs꿼��~iݽ�O����^)�?N*����b�]�7��ri�3�5�n�q�|�^[��fҞ��&�V�$���*�e1S��,i�M
������j�Ѭ��	��fv?u��A������^�a���!�[;��i��P�k2춤�ؕ�ޖ9�pD�L����aN]�l/K퉀���P�}=�5bs�E��iٮ�d3����u)�.�}a�PB�[2l����������U�tM��`���O|�F��� �C��,�� T�$(&�S�61�ɸ���e����x
ȏ?~y���޶���N�-�s�#���Ck_��� *|����=�`vհ���M�����r7�(ȗ�yi7x6^� ��[�1X�7:����2}�Xn�#�\�ö25�w�R�n�N�H3NT%s��e��wPP簩����-=�|FvLd�[v4���D-����)�X������_����j��偁A{�ҥKl� �D�g���o�t{���'[Ƚ��b���$�.�<�>�r���r���zaDw�nCο�y��/3�1�kL�/�,�Ĉ�7ν��|��9)���) �h�M������^w蔝q�87w�ސzͦ�p6[͆:�}y��?r"�#V�:zS�S\�+^���*�?��7�{w��<[}���7Y�I�xq��b?���r���'E]7�eT͒�����r��cg��j����& pܰ��h�0W�U	�Y5�m�'kX�I���Q�*I��I{Fg�D�p}�_
A����_�Zs�B���D��(L܀�!V'�G@�G	�"**�������pd���8L����K�ti�2�$WL1j���.�b�0��
%��A�"&\�x_T�����\�z���?ٴG�4�]U���= �.���dڛ��yVS��q]��]�٫�D)��iCV�S}նQ�e�Th�xGo�.}�HmO���&�`��ȯ���*��Az�1�|:�HS:X�^�1������(b���`�1�).R�l\�l��d�%��I��w��\���,Bij0��X�$&l����?�d����d�T)Y<zB�������p�T�7W���l,��VDb�^8�Adm��ы���9���Ȓ2)G~�1l~!p�o<L�O}� c=V8s�h`ܴ��
=`A��7��껫Ry�>} i�|E&|����OM p.44�Ƭ>@�ֆʒ�(��aXo��P��7�� �j��
=�Y甑�W����(�����6�D_�M_�*(yO\����erm�0��84H���v��rqj$C�y��R�R��ҩoKA�s ݌��F����ux�\�L-!l��jʮ-x��_��b�� �����
���}�F'��dK��e����k�;Y����X\�$��>^y$��۲��)u��+���<���V�F~�٣�Gc���!�+#wrc�T������� �X�鶺���K�[y�������l��j��H�Ci�q)�:-X;�(�?Ԥ@�G���V�@�hm�u���>���m��?B2?L�}��{w�&E�P�c�����KY3B�
8�[׮��qO	�߷�Hk��vsO�}�ֳ�2,�f��v��VNн��״�{�Z�iݫȰQ~Ϩ#+��)Z��L�̒$��]s �X,�N���j �S�ﰥ�xR�ݙ��5-���r�Ϊ��!�k5k2����FlGl��y�hفM8^�v����q���X�Sܔn��Q�NW��	��h�k�c�g��+*Q�� #iS��p����Q�6�kc�'�"�ޱ���E�
��y	8Qg�p��MT��~����=�N�o�.V9��A١e�ɂ 2H�����`?��� VTYm�{�b�645}�F6	V]g�}�p�.����C>E�$��'�ײǵ�@��rm���(�e������*ILqA�Lғ�7���*l�'ʜ�mh����d%��-<+L��Hɑ��+���e�x�}�8)�?��l鳯2\�v���J�a�G5�9$����6�^�!��~M�O$P	�V�x��y�� �(X�v3똪����� :��	&�w�"y.>"Á��IKh#��n�jy����x[�[H=�BqB�x�A0H��,�ts71��2 "�f�4������k�gMMVY�냻��A�8�Ahs��H�C��ป����������ʗZ��;N���SP�{�L�K,��CltT
��He�� U��A�-�E6�h�+�r�f�Ղ:����[D=���L�m�P$�^g����*%BYq�k >�
"�۷o��mu}��ʨ�c#O�h0a �`O����zA͎�|�:�B1+#LS�<zbY�I�ʩ���S��>ͬ�{�ƿ0W��z��\���d#�wZ�EJ���R+�&�6Jqւ�|x��@���">��x3̘$S��-��IX~9��O��r�Kw�> ��y#�"ș�l#��3b��sSH�����1)��$��xB��%T�N_fU��͍f�'�c�M�3K*������s��e�����ﲝ��Wdan����;�=H���"�^>���zO+w�j��sg{;����w�KV��D)Z��C��@��*� �5u��\0g�¨;�!����Y� t[�rO��'�2V/h02����YH��p���ܷ���$:ФĀ�x�0|��Q�&�3רՙ� �����j2��s:)!d�ɓ!�	�ۀK �
�Y�
�Q�;��Ҫm��k �������17�Z�QG�LE�$�⚳z�UHr0AU*��?�	�L�m�V+�� P���kp�S�N���~&ph]��N<�������3�X�-mvQҎ��'�,�>�m��	N~�$��Xk���V���O���k�GF@;F�
���Y}�&�X�LH�4�'�~dm�ǂ 00=�!��m�.�+��k� �=��=�G������[m��?�2��@�9�<Z�7n�`�q��]�����L�AS�&� c�1[4h��2U�I�gL��_Р6G	���R�(ːQ��6k�2�=y��]R:P�]�wp��d9<�i2ޭ�z���r��m���?':����I�X����&��H�l�4k��kz}"�JJ��F�~Nw*D�����l<͌�N8��HzF"�<�S�#!ٙ�FQ�iXc4������.�|���b55��P%�$�������	QaOߧ�8ݬ���d��4���	e�u ��R��Xyszz���@ȚFN����*G��Rc.��DPҎS�%g  �����jߦ&�pIG
�����F�R�n`�yĩO�xA7!4DB�a��^�u��vdo]f������\�8�+a�ݱ����'�#-���.��ڦe#���0`��� c�D�m��F�!����S���4�,�#��RԘ���j��r�X����˩�Bzi}Ny��|ZU����]�����K�A-���p'��MG2�DؐR��Qn}#����y�D�0&!i�:�d��^SkoG}a�Q�`�O��F�`����M�Dx�a�^��}W��&MJ�6~�O�~7�0R�������R���2=���/d`r��sBp ���C����IC�c�U�U�� DI^/���`<��l��D��z�l�)K;3�3_OJ�e:���5�4��TI�A}���g@<�{���"��ho@ĳ��:�#��(���,VF�����X�@{��i�nHy�>���� ��F�������ԩs��`M��9 ������,�4D�*�
�7J�{��b4?�Y�)Z�|�������>i02ć@T�I-����-��3iS�q��7bT�H��S�׵�����!�5��i¡�3~�� >*����N�m	`qb���hk�S��J�iP�yr�C����V�*X?���.I�s\���133��"J����k�&���O[@�`I��)����Z}bN<Voqv�R"v�3Vo`�~U��ap��)�A{;��?<K8�#�0}���)uޏ>����f�A�fn�	�������ݼ~C�\c�Bf�l��=�bN����	>�l>��0�M9�?�vU���MNpZ���5��gf�2=3˩�W_����wo��k�m�UM���ϰPȸ�>Gڑ��^Yս��_o2pFm�*�et_��C�r�<z����g�_mN�ý>�@E#p� ��LJ[7QBJ� ��~���5tZ0�4ꩀ;ZE�B�Jw8W��nܪB=;���$v �=~v-�|&�F6E,P�UÂ�Ym˿��e`����5�K�2@��4�~y��|֮���Lj�X !�\&pZ*)3�7@�/b?3�d
�I�D��i�cWF�bĞh�1m�Ȁ�ԳA%Go,�o�L��c��r���u�C��H>�̓t^ԕ���� �B6�w#��,#ޫ�	����'h����m���E�4w���y�g��M��"��z5* ��~�H AΖ���!i����4w�0��,��2P'�B	uO���l��rILH:ÎL|9��lU�>��VC_C햴��r ��@��$�	CGe��8!�mzǚBCr�H����@�n��7�+Z{��ǘ4ā�����Q�F�Q	0-$�;G���"������_&0�*��B�K9;�k�5����ʁ$�J�=�Pb_R�8�I!-$yji�2�g8F	@(��A�AY��:NL�
�Z)�'��z� ����h�t�V�,��w���Zʵf�c�2��d��HU!`��GmgK�\������pV��̡�6��h�7LlE�ϕ�h��N#BI5�y�.	�5��T��Øc�q[����ʬMy ���ǔ�p`c���$F׉vjS@��x�	�Z�p�H����~I��l	t���lbW:�,�냃��^���Or0/2�߂�1f�}y��vml}���x�O��聴�Mğf�Cj����oTpP�O1�7�&�`~u�D���N����,��C����C"v��� K�m�C�
DU:6X/2P&4^4�~#�Pk
-CK�F�L�&�Y� d4��P�t�8u�۴��ҡ�.�t�/Y��I�� P�����w`�je�zNG��ɱc�efz�g%�~ ��A�7��,�����o�;�C�N��8��|1M����&�`����$TU�����y���^]}HZ��9y������"?}�e]�@ʕ)V��t2��γU���-&u��U��I��Q�ڈL�"�|I���\��烫�e{�)��ǟ3�\H��_��	T������Z�ҴO:=]�_^�H�k�J[+��]��d�1GSY=D�����aR�w��K�M�G�T2��H3���;��Ƞ쪛�;tk��,����8G���6 p0�������2�R &@ٿ3CҪB�B���X�������`���tC�he�&�n����2R/@ac����:�H�R&�����|�Fv�P��q�WZ0+�u����ѥ�do}MN?���d%/'�x���?�07~*��i#+  ��EF��0AN0j޹sW�y�g�}���tͺ��b�5*5�y$�jd*�Cs�`�2��W�be_ �
)TU���ߒ�|	��3T���G0@'�m{:R'�����}i�d�}�zϸ?�SO���4 H�3,ʼ��%e��E�ltF�%t�Ap3) B+,�ұ�e�}6��{:a��<+��{�
�.�A�Y;���@P �`��-�$#�bc��>%/�W��ޞ����|?>^΂� ݪu�=<�� �x+L�[6��G�O���Ah�0qƀ��������P�6Cq$���$�Gh&/\��=w�_݃MH@�l���c�6�6�� 6*vp��#^���Kd�1@��lB��s�����.lL*�E)�d�;9`?;=k�xF �u�E"*���x��]_�;?C�����a:}:�Q� �����&��S�ƺp��y9�"`Q�ֺ�=�����P��Q��Z�����a7ӷqZ��!�m��04[9bX0�Nk�^o뺃BB����Hx��\�v��:-���ܥH(��QA%�hgxT"�k [�j�B{��/@�!�;�F�n�8�@��l�+�=GJ�T��	ˌ�i#�=�������b~hy��Ա�Y���TY�i9�v���9i���aϳ�`�~a~N�[���<�
�J�sLK�[D����a���Vʕ(��6���#|Z1y��S;�MTq6k�֫����Z]�J�J��焀ZO�]�ޕM�qf67�5��k�X���ҵ�mN���������fO��~��\ӗ�Ɋ����G~������i�U���X�!��T�����D���㩩T��W'�n򁀟�3O�f����.�F��ۡ�(��AI���(�۴YyX����Ț� Z:�L؃��><�HnMAxHʅ2�[P���F�-���4�MR�h�Ӎ`r���@���YOU�@�� X���$��֭SsR�Қ:;�52@g��V^���QJf4�6�t�x����|�.��_�u;#B�C��O�k���L��ict$p�#�������<�ا䕗L�Q�0��	��|���/}A��F%=j�!堠����mtp�`���ȡ9�Y��(�S�0� [���l������Rh��?`��6�~F���>���a�Hɀ�4��3+3�+�?)	�i�-��f��% �ĄO������,Տ�aJ��V��{�����-��8���4n_���b�Y<*~�r�nh��Y@��s���r�%����x��qe��_�:�����񩤂��[�scz�ئ$ �1{���չQ4nƬ�^�D$�3�K"�@� 	H�gR�� c\�7�qϽP�`\r���?O�\1�X�ŧ��b�q4��R��T��Ŏ�4Nμc'M��s����G�Hq9����0D�I ��P?kd�L��y"*�&� 	p���O[>y�(=Gmܣ����&��r����V���č�ʚu�����#��ϩ'������=�x̶�r�`�W`&U�ĥS9�qmS�I͔�.l�}���`�YL��c�u� ��רׄ�)���l��p{�#/���A�I��[�b��AVa�zmݞtۚ,�i{P��^�%�06���3@��d	8~�I���gR�U��E�U6�I�h�L��6���e9<7˪1>kvz����ɪ=|�Dk�/�/��.�������g���v\0*�&�*�;��z�� �\.[0��N���3����7�x�{0�.���I����YX+H; �>??/������p5�벯�,F�w���V�U�8\����Kxŗ���y�'qҌ|^!+hd�.��� �����o�B�S����ܼ��[��WqF��&��7��A,�X<u��`l���_�H����d�{����f���������ˑ�e�}pK�>�,�Jk/��M4>.ӝr�f�Mlֳ�5�?ԁ�Pw4�i�Y?��iY\8����@���^)�ӓJ	��
7�k�3^�xI�o[�e���:u�#�Wۑ~'G �8(Gܟ�Hڵ�׈��*஀|����S)��'�1r-�ȷ5 Z��!^���9�~G=y�<��i�Q����ȹ�.��;@1r�t�Ѓ �O[���j��	���}�ꗿ"/��E�V�c��%^g�ӐH��e^آA�ݡ�C����wXR����.�SpA �E	�"t��q 84�=)�G&�x���!	�"N�Rh�,�@Ȟw�h�'�mj&v`YB��蟑���t���P	�4�	�K�~������!�ȡ�)y�ϓϣ�yWzu5���u����1'���$��ŎҞ��y}<WI�sn���'�V��E,v�xGL֞/�%�^I��$!	���5�W�o�ƕ
~n�oc��=S_��xT�.�Ǳ@L��/H�{.�}�%d���TBY}<���a��7e~���[xX�Sq�⏽�U�l�E��`�(N1�����5.�L�a�TX��~��,��&'�R���~e�y��ABx�R;r:W�8l$b�;�A�] 
@���ɯܿ�Vl���S�Z�x� ��"4P�����"Q��4pW�Qȗ��{c����^w7�>�ddc����L��&�M�I�;FZ�6�w8D�W��I!�O��eE�j30�R�j���#Py�&����hs�i�@�w����Ge�A�O:5�.��ȴ���4���iM
���/�C�j��:=3AE�V�!��[t�U���&�ط����YX��8�������ٙy���i�N���r�"%�
ԡ�z�}�0�*9��,G�Gr��GĶ̫O:~�>ڨ�FW/.�P�f�;��O��/|�K�ՠ���V����C"K`�(:�(��i���6���r���Ll�zm)�E����Y����!��s`��f�����?Ib���Y)��R��e��&�"�1��G�A���ɨ'kd{��z���Q�*1}��D�E���렶OPT���`:#�2~3,xž3$d�5��h�������9����GyP��D��DK����������Y�>"�}�i����YѠV�|�]������n��O=)����BV�r��GN�������~�����o��r�iqQ��/��~�J����_��O���Ȓ4y�n䯿�y�՟�!(��}F~�k_�C�Һc�5��C��o��_��W�2����[,[w�bw[��F�E���#��z���/��i��N�{�J��/t�h�؈�8砐�㰟<�,���!�#^�u�P��� @��*6LB/�2�πh1������1�M��<^)m�Tt�����=�+�Ap1h�5����C+�'�B)�au�ҩ��\���8�X`� ȵ��~��9�8#��[f��,�f�n|$�:�J7�=s8|�n���%r�$Í�l�MؐU�\�`T�?��;�Q"���&���ص�a���P��M<yI��̐L�6�����bd�p(��(��/6ن�c'P�{�#�@�W;�m|�ݏb���z�S��5�q!��������߁�(Y-~-�Fh����k����$47�N���^����z�@�L���U�$1���3�y�|Ķc\��84v-�ȵ��d��%ց_Ã�o�,�S@�C�&��p�m�Zq�����Ud\�1rk�����.��\�#c2��׋��~�,�`���h�a�0�s�:G������hP�ܕ���=)�F佁mÄ&v��Y�����v_���F~N2�D!Z; _�&�t��m�K_.O0��Tۭ[��Fah�?� [&��g>�����N��/��(��<55I��cǖ8��	ɶM��a�So�	GN�Ǳ�[��s�rKG���SB�{�y�������,.�������Ǝ|�?bИ��A�c�����\�TŒM�	TTz�oIn{G޿4d2I	h���A
�$*0k�PHNm[��L&�hE�5���1^�������m�T�vf92���?2f�t�0J�s��_�[e�T�ĳU�G�E���e���y̰c罥s� ˘���
ʯ��A��. QO�yD���e�������g3���a�F�zhbu����/�)y��%y�'?���<��/�?��Զ�套_&������>\��~���ך�7~��/R�W(�n���O�}H>��)�r�ĚIܿtX�}�QN���˲������g>-��_|U��m�y�|��O˴:����ˍ[7>~�� ��`YO�xi�N�&���]I�pg�@ՉrQ7�#��?�Yj:��6����f!�/�Ц[��b�ϑ���2�>��o��t-oʵk7���� Bh9��@÷���� ���.<�,�@ �3���b�~A��� f�3�>G�3,�{�F*�+#á��5	��_�|%5>�O��VWn�]3�ϰ���fmOn^�����Ghz��� �Z�{gd�M$PW�h�(�1o�xcÏ��=���Qt��|��4���������_�����@ptPy Q��iW	�|:Vֻ\�B�� +#U@��*�8ę��օ�\U&�%�@�w�����{K��H㶖[� 㯃.@l�7�L�3��b\������3n���=n�Zl����6�x��q�L��%ϰQ���8E8�B���Ӈ�&���b��N�����|���=��>��IPBs�T'�wҜ�6�h0�8�!������&�lB�N��WcW�Y��Ve�ViZ�����c=$5u�dQ%N�+�־LLUd���ŮT��L�B*E�ݒ��<���ϛ�^�H5q�P��n{�����L�T�o��ҍiEeD��74.ɡ�K�9EyHR�I�ٙI��Z���ɪ~_�v摇�'w*�H��V�����ϑ��Ydg ��}'���$�$5�TOma[�F�F�?5#�=v�T�� ;4�I������ΰr�*��Ϋ�3l�&�%���&��2RL
�� շў�|N��]E��G]��!�]��{���y��C@���� ����6��ݰ��P��{K����O��V�6�A�'J297/��S���ש1 f�5t=o{�����ik����
�=��Q�
��4F��8?�R���]���h�7VV�}`#,�#{졓U�����+	��bT3����S�#�>|Z���o�!rs�|�ߐ�wV��ÆE��?��_�G8!�w�S���S��˼t�]��{�i)�EΟ;'�y�$��n�H>��g��Yټu�%Ү����]=pkr��%����5[�N̰z �799F})OV���<#�g�����f'�D�����<���l��A�t.⧁3�op�P�CZ	���s,	?��Y��������?3H�X3�@�@���*!��x֒�aEV�V����Г�)�����L�!�ĉ��~0��b�7*ёQ���.�0s3U��(y+r��)5�i͈����ݫ^�z��kdd_��w��?��9=��{��:B�	����|8�ĉ�x�J��L�$�A\��d�)�Z;��@-�Atv���1��L�d���=��~�{�Jd�8�&�{ޗn52�IB�N�y��PUC�p�*n�j+g<���$pm������Ecׂ��X��?	�l���wSE���x��?�c�1[?��>4�=�0�I�ak�����e��w�s�V�q�$�'�H�	kW�w­ª����� 2��Q�]"	<מu��q�Y�6?�m���_l2&a^���W��o�r�<k]��>��CE qh�I�cjܛ�+����a�#N;��,�wn˷��]YY�m�N�C����)��R���<S���fei��IYJ��'�@8n+űU�A(=P�#
�d2��Nc �������-�{��ѠEmI�+s:������G{������΁��Q�Q�'dE�R,Hs_̉�:h#�k5�8�>;7�[ǿ�u���6�Z�+0��:�,H�)ؚ�KE�d���W�ay�()'P�F���*�&������_�Y]ߔ���3s"'N�ⓄF	M�0݊
�Ɲar�ł�zU`i��sD*lQ���V6�.A \˨��6����x�^6�ǲ�wQ�����.���V�r�Y��d>~��_�H���^Om>����}'�ӈ/��Wnɝ[79���
����PB'�J��8�Eɋ\�Ϳ����ʁ��h�l��~m[�Ey�чe����ڦܺ�"7o�у��`&���	��������q��Ǫ��A�LZ5�kw�`L�?�	��wVd�9������`!���OKS����U����3!]�@6u3��=���呅i�����ޓ�ߐ?��?���-�r��\��.��_n�kƓ*�GI׏h㏂i'�FP���>�q�/|�y���=Ҩz%�R� ��S��X�͸j2j�]fsɆ���X��7����}O.�?/Y����ϔ�$��Z�����x�o�jK��̹0��ǤY�.�!�WP���x-&>�q�"q��(��fb���P��3l�0E��
5��8x*�5�P
F6���NNO���C�'ZO��>�PS@΄X��;�hh�1���&A"RGn�$	�}#��(e4���G������lp�:d ���I��m�z%��a�k�$Z-F^�V��o°�6Ř�ap|K�&�#I;9��pX#�\%q±�b��%�S�M��Ԛ�x�q���8#�&��ʪG���}G�f��%I�7nq�T���9G�"�����Hn:k��a 76������tO关=|O'�a7lD����X.�����dm\��_s-{8>��h����Zr�wLl�ީt���82�g��2^O����SJ�� +���o/��%J$\�|��6����RԬ���c2�6ty�(�g4i�gɅ����8��e4���0��>�ݺ�t}*��qh��U�Jo${}O��=	AЦ����)�^C
9u������nT�4y^�[�C󳲻�)5z9,e(b�v3h����?Ɔ��=?�2�^��Ӈ��`=0�}�}_ d�'�g'�"�t�|�y����;�>Z:�([ۻ<��b���"���su�����]V�u�g�ZQ9��?��Y��K?�+z���Ϡ�@�r�-͐2�E��:�NCU���VӪ�<	"+Uik�� �Uʡ���u��qaT`��ÖLNU9%�U�t�\���>p�r� �)
D;' �ؕ�����'��l����	��\�0�e��f� \�H���~M�8s�ɳ�}Z��ܧu�ܑo���ɤ�Dbkg[3����=� ��P+�hQ鳗>8�����p�e&�]� �?}VN�<%ǖ��PT����9�̊Ų+����PQ!��{1��������R `Z�[�����s�df���?���rE�|��(v(^� �MV <�)���eo8����3V["�<%#�I<��?�{�j�YN>�z@��_���>++�n�`�<�^�o-�O*�=A�0�!����q��&�gc�> fJ������5O�qdzpz+���m�'����Y�>x���y*g����<�MA�����yC�}rfZ�w��Ȋ��bZ0� �̱&={�l��A�p2� ����	 ��`�	I�l�8�%�#z	pIU�솅�A�Or.�Ύ,�)W�t�KL�fTb�1g��ȷ�]]L������Iԗ��J���R|q��kiËg%�a6�'@c���}������*���D�*���tRm\C*02���2�I�`���j�`�l�y@_���t�3I7�7>���E�T�8g�fy�� 5�h�'-C�q�"�B��bYEtU�q�G�Ӄ�w��\�od���A��Q���zU8� �c_�w,���	l+��UV����i�{�����mo�}�}2邆 
'*r|6/�K�,Ur2��K���E~fpz�`�VY�i�a$$c�(�gc����]��lY�h9�Qlv ������m�Nm�Q�{t�X��D��T�y�}LOVeQ�oW~{wG�_�a���@*j+ �ET�f����ղG��tڂ6�T$ ��	lǂ�IQm���jOa}�'���)�Pc����%�����Z�����O�g�g��������/�m\)�� 9}��|����NU42M2�I�5��C�*�Ì(���$�������>�nl޽!�;ui����bgU�&�}�u�>�@�\��b�����l)'�{W>�zY2�3Wf��?���Ƚ 6O�p��q>��J�R�+L挚C	� �b<��OM�^�*��?�x�a�x��Oə3g屳gȴ
���ߒo��, ,k4[����®�����$S=�dJ���l�/J�`j޻|E>����O��N݋��}���祧l�X��}9�4-��$����=�x�!p#]�f���~ ��ۿ���������-yࡇ5�?"/~��l��zpA�����Wu�����x�ᇜ�EZ��O�,T�1{��(�o��a2^2Zf3����ƕ����yy��'���N����l!K ]�<"1���^���$ъ��@������Li��E6���SAZ��L�*�s�͉s��'��N�dyT��N<�Y�0ڔ⍛r��syr��t��mT�`P|�\�����=��JC>�S!k��=`��X0�ޜށ� �`��}���G�܀B� �q��SIt�t��8��V_�t8��9��v��W�f�<4e�4�}�R"85����Y����[������()��u�䌾8��l*cZO�{Ĥ��L�2�o��N,/���dtj8��0�(gc�����$��(W��q"cOd�A��9)�j�gbAT�`�m�Jk��8jq,��T� ���~V�#��d5�?�d҉C�u.i�X���R$>�M'g��� ]��5� p�� �5R�Tb-�B��Ȕ1Uұ@�3/<c,8Hu`ϵq���3�:pe�6IԃA�{ȸD �+��2��&CXKd����Ɯ�=�,Hu��Z$�:(�Y�s��C�u_�)؃��W�7%]�#S92��#��L��Z�.Y|q_`��[�)��`��L��T�0X@L��Bh��:C���kڔtvrª��@�) ���[�n��{��H��g�j9�Y�=�����\�@�H���6u�g�,(F������mfn�Ո-�}�.���u�Q��y�&؞;�o���E�Ux��C��+��Z�p���,�M�deB/")�c�SF�s��U�yp�@��v|��YVB.-m�ܕ�)3Q�������14-M�iЇ=��ݷ&�85QA``���'�`+�<}�41���������Y��ptd؃��B��A�/TO�8��f�~*$'2������Y�� �ҁ?���8+'�g����ybT��h�Q�(6���˅�?��O����59���m���%y�3dm�v�%�=Pi�� Ϲ�5!sr���\��*�:{�3�?��y���K@�~{ o���<��	9��r��F�5�3O<#������_HirV~�7~C��Y�@������@^�٨w��a���-�!�]$G�2��h�Y�`�����^��e%g�N젤�Jȱ�i�5�w=T�Ok�����@f�i+�C�ؘ �9��E.�sO7�`�,	eYbQ ����+`����	Am`mA8�>�`0-��@�FM���W��_��)aؑ-��%�t���f�O1�(����Hf�h���q*H8��t@@�8�XI1��lG�{�$��M�z)=��*&�uҶ`˓�(`%W&�?�*)�IZ't��>M�F���{�����z�yO�,�5�c[���z�����uA��6�8i������_G	��Q8{}vXS�1�ʊBdU"Ts8���*D�К�k0���e�0�wV�Ԁ- �h��*T11����bI��.�Z��~>�P�DPG�� �{��t��� �ŵ1�z�pM-�s�p�1�F��F��g�J�1��׈�n��  ͤl@��
�&R�Ŭ֨�˔���A)�^mi�gf83[�)�E	�\ [F��VyC*��շB�@%s�����(�ghB�'�]��	��Ӡb�:����ᙍ�A��X�1�����h�{hm�MN���C����/�bY�~d)��U�|9ř�QY1
|��Xę ���`�&�$T�!a1꒴s���r�J��x٪�ewGZ�"QB���������α�B?��\��}xLOO2h����Z΂2�.iJ��x>h���	+tRM���5�Et݀�� ��v	)"(�1�V�5�4�'�f��p����yNN��0k�H%A����$��&�_�D##.�'u��o	�ɚ��9h�&��0[��=&'���W�� ��#LLO30�k"��68��emR?��(�.���D��N���!����@��޻#����$X������%A�0�I�9�CR *{�\Pf"8(��@�S ����?����jWn���?KV7k���ޔTiR������3����jr�-T�����|��ْ��&���B6�Ʉ
]�	�ڽP޾��<p���~�7�����tuR3Ҵܺ�-?y�<����{�����ӟ}��ܸ��II8�)��o>'�������@'쥟�&{�+��%5$���C��^�����~U#�+Bβ�A�*���x�ˋ��F���e<��J@³B���q�bm��S�ar��F,��������0#@���b��lW���<=�+p���<+�4�b,��2��A�2�@ �a���4���_�(�N_6��pb<�P���<&:� ��o��iL�4=?O��l��������ol���Q��9`����ս��2Dd��攐e��a�ZoG��g%�شk��¬T�Ɂ��1W���M�1�Ψn �A�>dy��̠-��)�ޘ�]`/<��Jd�`?Τ0!���A������
��_�hg䀷E5�|�`��Z�	�k�mA���b)��Ӏ����Ԅ��0Q "�z{O��%p�U���LH3�^� �`�اq����T�`����ֶ��Y�Ů�?����X�G��T0V!G���W;�j�^o�g8�s@j�O�YSn.Z�A�҄{��w�#b�s��h��+�k1d0��:��}�V�i|Ejg[�����)JQ��X�i��D���`���aLU���9��,���e�Y�bY��Um�F\���v��jl00P.����Ŝ$9�g��tޤJ���<)�?pD�VSRN���U��S���&$�f�J�ѠE��P���`�-S���Ī���T�6��>��@���� vR�;����p]����~�¹F���uYY]uA�H��s��p�5	����ɧ��۪�H�DE�~w�@]����A\��hl�p_��~O}���~oD"6`B(h�p�� ��f��7�c0�����܌h��������s���''8:���0�O���4���	}�1������9���Ӣ'�L�S�ܿ��*�� ��k��j�6v��A�1;�[oq4��S�5�벯�~l�sks�@7�ʳ1��o���J���	�a��F���߭�s�Wu�r�ȬL���(W�o��s�ڭM:��/^���@���/ɬF�^�"�����_\���oI���n��xInܺ�	d�-�&����EO7չ���&���A�#HR}w�K��![1#C-�YY� ��eF����^$�g)�>� %�q�k�ɏ_~E����uh���	퉜!���_ʲi��gq�a�Ӷ��5��y�*�/�U8J��I�>��g9)����2�L����z�x��fLd�[��G\-h��B���A�(�������g�Zh�S�#��s�����׀�Z���5����]���5R��؟z�A�ug��=G1f���|u��$��`ͅA[0�>�B�y�S�l�o�� V���	 �o@V�x��g��y���i�� ���/��w�DzP�gea����f�:������>�b��,��K�#>u��
<Y/m5��ʺ>�\��A�n�I��_�C��*��� �Ef���~]L% td���x�O�LN%Dd�H(���̝���{����r�|j�x6}U.�=R�e��ImBO�N!�'A_Z9�`+3ZF�Pd�����6v
��6^l�Ղ�Kd�|C�-�uޒ+K�P���hJeS�pN�l�4����<e'(ݠ�k�ɺ�"/�8*2h�}�`t@���`�z�M��p�I�zQ��!Q��Q�\a��dA^��[�K��{��2߻٨i5�s���&��jY}�,�!o���j�D�J[p�}��yƣ~�6��� 	$�6*����ײ��MN˼:�r�OiN����t>�K��b�D���T�7�9P2�q`��<S��R'N�V��i��~�Ɂ�u�����^M}PCJ�W��7�v�X�UJT��--�}�Ѩ?ރ	�� ����������4�g�I@�6��ow-�Bf�Y�YC��B�{�]��&Ɖ���	��kB�QD���> ��g��[YYa5���e����O���wF�ԩS�|J���B<�b���d�r�������Ӊi���%��Zi�����S��z����e[�v����!QhYNr�<h��c�G����h��6C�2!�Az��� ����;�rk�&%�1��S#�j��#�:t��8ݛ�{r�O����l.Ϳwj;��2zЋrgm[־��|��˂�SG5Kd�;�}�ޏ^%��F�B��J�_!�X~��E:�Ѝ�����s%�ՠ^�-���%:=!Tj�!h4�RA/2���V��T�z�i9������I���D�1b�������h���TR\u��qt/����vw�H����"�eq|�<�Ȃ�YQ\+�]�822�rZ5�K�=0S��4Q%�Տ4[��o��~�*M}v�����vG�f����D�ѣG�䩇(5��]�q���B��y9�lˏ~�#��\3�b�e�C�?)��B�v��)*N_��Cʴ����3X�ײ��#�M���2���Y�+-(A���t�1�:�VK� ?pSL���{d�է����Y��T�����
��e�FJ��j�5�\F��g��K\��:�@�Y��s�eg�� ҹx��OW��ݤ  ��?�gAl�R%.=q�|P�OA�[&�ٜfn�^�Y<z�8���3��%���$[n�L��e`槇\/(<�^  D~Ȋ��z���Z,q��	�@����V�R�:�k���!X��]�{�i��@�k>tT�]��E�ȗ5�S�I�|��$���}�Y94U��������^ ��N���E��g���-�ڐ�~�ܑe�`���壋����ՠzE>��!��Qaɦ�J�A�
`#V76նtYm
t�B�b}(��y�s_���<,}�K�`vw���c|�QQ�s��'�������y]s�n�ܾ� �����Q	�=ɤ�YN�Y%
�<�Q�us�.��~��j���t������C|J^x�|Ig �}��YI���c������A�@��k�4	��a�7��`�vpjr�U;�D�������)���g�r�Ċ��4{�a+��a M{`��dq A���LHwH��۷oK{�&��ot���J1H��
:�uja+z>[j�QeD�̽1U�G��ݎ�
FG�r�f���� ,�U��=���)4H��0ըIHJ� �vK��	��yD
��}Nj����G^Ə�@�O���*�b1��le�C?�F�x<�lo�H*��x;%[~2�iQrB���L�t���F�;�08����1�^��@��"2�ك?҄)ǒ�O�
� T�A@:S&`�݋���X7I����89��P���cgw���$����D��2��݈�M:!z�REN`S��e��,q��:4��<+��g�"�`���z3�1���4��QR=bV��b�0����� ��b�c��a����hXux�_>��ME��~0����f(�i�c����pz�����G���Ju��W��1_�ob
����4��kˮ�p���Ӿ<q�I���9��pz2PǴ���[��������;�dsLT��Ҫ�h��򩧞��@��s��eY[[�:(�2&?kL�9����)p�5U��n�*/&��PF��Iem3�B�VJ�2�H���MʪN=�/(i�]T*�1�	5껜�@pa�-O�<+a�&�^h� �N�b5 ̻ �:u�	��Zg�� S5�#�ܕ�y��°:���~�o�P/��B�"�g	�=��̫c,���tu�;`�p���%}��l�Z���C�k3(��� �;��,9���s�4�
��j[�*����]�"�B�{��< )��+��'��d�}Sv77X}�s8rK3iLhL��C���%�vO3�2G[��"�E�T��o�˯�W��yY���ڇ�d}}]��^���g����_��^}M����Odm5M���C�K�ʤ����TM�-ȓ�zF^x��rg��|�����!��&ԍ�| !j��٬ݔ���o���@zT ����]Z:F��죾̨�/�0��֘�=L�mm��S�&NC�-Բ��!ք�8)��2��d\��U�*��QT�@O9��K��O��(7��>��q̈cŵ�J���9�<��U�!��i�VTZ�Q����g4(���d��amt�JE��!�����%�QMK ���Y�qzqK��&��\#�Hl�y�X��L`w�{��@Tכ���59B���I�H��z�� H7
&�����`�L� ���5Y`c�X�i��>�I耾1p��Xw�2��66hs0%�$C}������׽��d�-�.H.���B�[4=9��9�`׍�d�y�`*����*�7��R^4������Y6Jͺq�P�Q��Q��h�b��K�нcmL���ѯ��x!�0a��d���� �ȴ��#��h�����O��x�=0_ay�* ���ǈ�P�0��M��C��{n�(Θ(b��3z�F������F�ý3J
�E)�m7=�ݡN9���������@?=	$�6�J�LI�P)��?���,nfa��a2Ox	C�#m�{^�B���D{&��"b@����#�Ν����Y!��?(߲T���o:.&"�Rr(&�b��`q�1���� �z�5#OG�Y8P���މ4P�1�
!H�F�СC����z{�}�R�D���\Vg���U���F=_��}���M��S�?E���N������ɀcw�euuU�e_��p��=nX^���!�jV��h@6����10(h��-��~���AI�@,@E�^���dU?��<���nߺ&m5���v�C|l?F��5K����}ԋ�
�L�TV�48zR�����Z�#���7��x�c����X<r�U�������oq��R�tL~��j�O=�4���}��z��+?��u�楫���Ĕ|t����^Ǆ\p�iX7"���8qR�x������4�ma����j�]٪���9����##�C@��mB�����wQ�FQ��]]���+�Y�B�5?��{K��:wu��B��9�]�!9�vvk�q����>.�gf�wޑ��ǐю}���g���MV��a�x���>�6Q�Pg�����7ސ���8E��f5
�z�s]�D�z��j��*��Sl�@�v`�kRÛ7�IY��l�b��LY��,��ex��1C��NG,�0�X�al��w	!$��FsJCٷ���l�ۺ�#��k��/Р ��~t��~���v	"����p���s�#�q�j[;TSc>���=�6��u��^L���ү�s�-=�yv5@������ށF�����j7��p���hx�Ʉ*[Z�&-ׄ�*�3h�*a#�1d������&tH(��-o$�0��*B_6����u^����,��� @�CV` ��gᚒi�Z��kc�G�'�ȋ�������*XmQ��ٖi==~F?���W��d��=��6kr]��\*��^��3��ţ�kIz��z���@�CHv�hH5O85�8D$��0!�����Ī������mD����i�=pS3pݶ�[���Sղ�9�ZQ�E=>l
d��wo$Wz]���^YY{a+�K��D7z�f��\�"EQ�DMhd�(y4r����d�7�Ȟ�R҈�D�"E�H6�zA7�}-l��Bj�̬�3�{��|_��#��@��|������{�=�y<0\�!,�쭃 ��-YF������82�x����*�X>�^Gw6�j T�X���:��7wO
+e��Q���!��1��8`P�����5Ւ��83&�E���D39�j��.�ng;�z4欶����>�c�q |H����/ ���!���	2YW�~6%�1��2\!G??�g���f�ؒ8F�# �� |/ʪ��
�#�:MIz
:[!�H�apL��J�/e�'�j��Ƹ!Q'nt"4K���!�-k�齏`X���&��-���@�zz���m$q�%�#�}CК���^��u���ǆ7r��t��L/���yh�Vٰy�\�t��`�Z#�� ��+1z�4	�p�^�۰�%���/K�gP�\�)
VX·M����@7�T$��7��R�o�o���^������� 	F�����K�D4xA(��=ݕ�=�їG���S��<��ݧ�/ KA3Ch���"�dv�ȩ�Z6�iM��������
d��G��iP؊�H��J�NP�C��Qg=xP%�(@@���)"�ܮ�*�V�&oM����ӃUO ڒ�ކ�����
� L�����8�=�Ad�/��$]��)��oD���v#��+��MP@M��JNM��h����MQŦf�s
d�nM��>��� ����i�ڛ����Gϱ�H���Q=�\����,������Ө�s��z��/+��q��C��K��+��
��Y��&`:'f���E}�\�[ݺ���Tc�M_'�Ih6?�q)���1�����3���A�*Ԣ��w5l��V'Y"F�HZ���ɿ@�P��@l�2S^�}�4�Gd5.����mt=�4�;�|�D�
 H��q~n�dWЬh\/��4�����!}�iV� ����P��Y�G���[L油-�;��{� �4�p9�k�p{r���#z��
RK
���De�����رZ��뉝 ���GV2�Z�� pt���ACg�#\�F�ѡ�Z6����ڵk@t#P�*�C���zO��SP��u��W��D�S���@4m0~FQMpBIM��nOI�ִ��@���9�������O��]�����^�.����=��'@�s*���V�V� "���f��~ˑ��O7+��*�n*}XJP0���DY] ����H�pJ"�Q��K�SF�#Zh˚�'4X7M�}Hl��n܄"�$�3�HA�'�r~�S��+̨�]����`�)�+t!�m=��0� �'��!��]p^��r��ʂY�}����0 ��`��v��0	Ӏ�E���
2 ϸ��z��� /�h��e$�=�Y�f��TW��ѣ�~ðlݵ�UN�8�+��*�/�1
������i�&�\J�O��e�qs����z0�0�x��� �5L�ԸY��n��J�BW 3�A7����2z3�(���2_a-.=]��48E��xm�B�ਢ�qA�cI�s�eƼ����3y���MM�ɶ]�ɫ���\�� �լ
����M�^���62�e9�d�]�r�Y'T��QZEyv�昌��Ԭ|37z��٩gX�!���������.@Zm�&�b�tk�u�EU�������1�����@u��d	6�eIf43���~��k�S�Zm�|=��X�F?ze��A{3 �ס�t�ۄ6��:���<y��)�E⚝E�������E9~�֖��ϳ��)���
�����~�Rqc�G]=�dvzB._���RAНIj�t�wA﹛̓P
/�\� �qI~U�)�����:�l�a��Z�g���"!���l����9fD���`j������X\(�����РV|]P~O�g�h�Q��ѧ�?���A��zp��tI��9�@p<z8��λҧ`d���C(V��_xG?�yG�f�����s��<0۫�<,�D��B]��a ].��3���.۫@�_�ٜ��K/I:�8z�g��YMRs��h�+z���b�����\���E:c}�=iu�I��bߘ�E�¯Xϧp5X���*F���?���1�|'��*8�d�C�B�@���z0�{nyyN��#��i`�@u�г���)krV�}5����,�)4q�jR��K��O���QBV��
��Qw]ewf��KhoV%�L����ٷm�*�Q#XWPZZ.�rМ��t*��D�ɤ�=��B+@�a��4QPlQ����0K ��PjҀ?�иߠ'@��.U���|�W($� �&>������L�=$�����p�/\�L�uO��aTO|��C�E�xq~A�1ժ���U]G��f�eeiY���׽�������۶LLߑn:*g���
����/��ތ'�� J���l`b�w��.ϸ����ɬ$AOΎ�bL$�mE�:c�������a�^�d�hbe�Q8� ѡgN7���J1v��\J�>�h���.����C�2=��ݦQ�t�$�
�\܀�\X������T0�N�FǸ�b��B_�meA�����'��q����3'0JڜA[*�j�{��2�����nY^���~���E9��G�)fɷ���,�y���O�Hw�bRS�d�"և	�|QYZ����zSLNͰ�x��}�v��#W�\��fp�l��e*E!5�#Pm��/+*�8@�lcU����C��Հj��|L�=ѱ�i#LE M��:=0S���3�8u��u-�l�&���)&�Q���e�r�k&<��' "�J�aڤ�]~�8�"��X��|/˵�'��e��9���C����XyCfM[y�|�=�U+z�H�j M��`=,.ͳ?�2x.�8��^�@�R�[yg�c�y^��*��yq͢��짣?αd͸��1#FX�k��Ơ�O�D�Dk�����p`���z��˃��,/h��v	Ź�����>d���Y�}۶r���P�xB[d���kC�􂼙lw����?��µ��O�Jz?b��nW�3Ƀ�\����vd�5�h?�r�Ua:�BA�žl⁃�(���/��'l�N�J|4Z����H��zaǦ�x@��] Ȉ��o`X�犼q��0�k�՞^���̾Q�K�����ʬ�
 ����㶕R`.�@+��cJ����	�W=�wMFv�*BF(1��Ek�
q>���t��1�QM�}�֨K��	�]]i>�/$��a�y�����B� o,��#U�V�؊w];��Pj���*^_��ŋ�
5II���$�z6ª�c��[���N2x�.����wK�?ZaL�DE3{G�>ϔZ���e^S��BMדƨl���C˘$]\.��I����u�l۹�S/h�l�D��4��MR�J2?_��;ST�����$>bEh	ڈ�P��&�$���>[h(���Uu�r��@x-�>�"���8'��QDE�J�ז�\.�+A�U�ڐB�,�����ڱ��1�-�-���(@�zs\���rY���K�)��
(�"�+hE�x�$�	��ɞ�,[uը&�ˋ�TqK5�*��i�U�����-YR������Jg�,�v�H��QQ	$����'�*b�ά�|L��5�h:U ��xXêpZ�������A�s3�T�v�ꌳ'Nۺ��ʈ9e5AT�D�$m64���i�ӝ�'�+�O����SׅPo�Y.�R�a��¦�)�6�e����[s[)B���w��5�h���L�r ��G��#��m`dё���}X��IG#�"�5E�"�,�4s�ܸqC�H^|�y�W=3�h>�����PB�*EBV:D�� ��;�6��M���1A�R#�%�ظ�|�y�{���Z7FV<$��8��r],ø�-	�VZ>�x;&q�J�
��Mq4���u6ErC4+5x�S-E�}ҭY���1�x砤O�� �4ΟQs�!8U��2�$[	شl���Ƀ>(ݺ��nܤ}:�����n�5�60���K*��g�V��Ͻ(���'��^>ל�����g����?@�����?���鷆� a�缂)��&S�	pbK�1�Y��Fz�r��9���Z���R���y�A*��H~źiيF.Kz����]�V�ĀK�:��?��G9E���Y=<d��Q����C�a7�=���ޕd���z���-�3��(��+�Ɣ�� ����F(�c&	��$��p�mꡎvR�=�$�������!I�T�U�XZ*u�ڣ�F���~>��A�����yVy|�Ө��ô^�f���Q��v|fAr}C�=!�Cx�u����/ʃ��I������Bv���И"����,LW�G��·]���8 3�sR(U9R�����M[슅e��D�������i���2�9	� "0i =99)۶na%�R\�f#е���r��3)
��tO���z �P����D[B����k�V�s՗�3�&�r�y���JA늤��{q	:Uʾ��d1����0���I�E�(o����c��0����$�����ϊ�9M�0*E}���6�Ju�r!ܘ ��>7��`_�����y��V��0�~�����Dao�{
���ׯu��>iO5	������,Q3` 1�X$X���(_�$��mCW���s�2.xB �A%`��	r�𞺲��b�� ��T%���/� Ey�O��{��������w����	��i�I�pM-hG���L���6&�t�t=��3�n�szm83���ݚ�

���n�b���uO�J
T�;G�5K�����܎+��ُ�cr�P:�u� �i�T�W������|�l�����P�@��2~�g����.�T.��p@tl}����&�)���%dۖu��{u�Uev���A`! ��v�S(1�$
g�c�y	�ڢ�������XB	�n�Cb��t|P��	�[h*:���װ�hd�s�Z�_q�,z��z@g�bzh�ȉ��Z/���.�8��m����T��<[P��[썢U���� w���t�ޱc���؄|�ӟ&����E�h�`CRq�3�	ׅ�8&�-�F`�M��B���z�
z8�e=@��֍�R�5'������g���Ή�ed�nyx�3rC3��Wt�7����s��=�i����,Z���<(�^'[��`��G�>�t�S9�.\�^";�n�/L˺�y�6un���3| ���K/J�Р��y�H�z�s��U��oʧ>�I��QFˢ�Y�֯_��X����lo�REM˄���@�`�Ϳ���Ư}U֎l�3�Oj�)*����uD$���Y�U�]S��A�#�C���c�&���ڴ�_�sRZ����1ن�5d�8��{�x8�\3Ʈ��Z.��������|�S���>�_��2?7���"�F��EU��	����xm�.L&Dh� ���FU�_�ȩ��zB�׌�5����1�#]��,�aU��e���R��	j �QR'�1ה�;ӲT(�?��3y�����IB�ͯw�6�[ ��?��A�
̮�{� -�#�R��֬�gj���iT?��>Y	c���P^�!Wo8��i�]�q�+HhA�I���𲂜KW����?��?�lٶK�n�$7&�����B� 7��0"}k�q4�ϴR+s���{[�ͩ3���mU�38���<��'8U4�7�#O?��lܴ���H"9�[��*�G�7q���7�'����F�j`jJe�i3�	.l�{�ݼ̈́$�6e �ɺ��l�������q���C�Gb�����.A\ULnV�C�j�X��2�����Ƭ��u�� tp� ��/S^��������cu1z#Y]� -�y p��{o��a
b�^�r�(Z�Z�!�ld�,���Y
�@eP�mY�еk�Gϲ�g֋�tRM�'��u�n�z�UTl�/����5�)��26-��Έ1�;�ќ�5L�l �º�"�+`��x�l�G�5
4���Մ� ��V��O�<iL�a��ޚ&�k֓��"����g��Gtd��uLP�:�E�I����%$����L���7A�圐Q�"?�� ��h�`�Ī�F=�L���,��]%�pL��j�//�xP��2������DQ3w/���n���X��^40�k'0p��%H�m���0��2��m*��)e��W�l�ZWqVF�R`e]*1bt�-�_z0ȩ?;�ࡢ@՞�'N�G����Q2�CkV&V�=qd�h�1���>���<���,u��Bi�S��fY�زe3��b�Q	F�_8����Ȳ��M����Md�[�T�s@sƋ7$?�NךLh֍�xL�j]��C�7ɣO�(��������Ĳ��t�k���$ʝ ��v<�bk�J�p]T���xٹk7�5 ��rk욜>{��jx*��,Ї�%����c��2sۣ�ޖ���D�KF43���*����#�?���/1��;�G����>n C��vݿW�y-��#J�x����P�$Ǐ��7�����!�=���͉I�롅�#��MM�hPY'�����a!=d�X{�	���=qKN�8&ϝ�Q�.QU���
֒�y��zK����]��˟��i�ڌ�����q�:����=*���Ə�F[3<�Qˢ�L���Ƨdמ��O>�jW�� GQ���+����{�ʥsg9Er��9
�����l=�y'�{e\�H��<���o�,WZ� � c��35-o��S��e�Μ|p��<�أ!s�Ej�蚺:~���?��<�ȣ�R�������?�֛��[o�=���>:B����D�,�s��Q�r����O�,��k4���f�F�3(���=z���>�q���qcb������/}�+�A�i&y�+���i���u��|���dҀ����=����O+@�{�OȂhO>��<���``�P�ڕ�
�p*����fܙc��2��J
]ZL���t礸4+�ZE�G|�#�%�2[��۪ɢ�)M����y�O��K�;�8���Ġ��<�X,����ks�%�����F�z@��3�@H� ������w&RY
�%��-�BR�g���g�^y�goe,/Ĝ��{��B��3��J������7�����!$��6D���U#v,��n���g2�g�=�[G-T�(&oO��70�]��z�Zl����H���~�P,�Z����-9|��TrB���}X���w�8U�Qp$0�|�K���P��F�h��$8�l��
Ќ ,gtm��v;�gi��랍N�1^���q$�̼gN{�ʔ�Ƭ�i�$��L5�����5������J���3����58��!�D��\([b�"i���b�c����JK��x�^L����XUs):c�5�b��@G��%`+�����������	׆��3H��x�Xu^�h�tL�h�, 2��E�/,[G�\S]I)��0��~���F�h��ķ�߬�D0z����;wf�@<.��0��(�]A(�4�����]�^~�����iA1M���m4f�jKEfI냎S<Z?��� 6ܟ5 Lt�=��3�md�|�Ͽ!�7�J���ź�{321_��E�{Y�x}L�Y�=GV�A�xho���@��쉭1�	�,����G?�5k����@w�5����R 03�=�E���o���e4�![�ae��Z�NW��~�#f��[�$w9q�q������%�}�`���v�&���1�}��EA[E����̝y����x���4*�/^!`�_M<�B 	uT_��̅�ԥ�d�خC@Ey�W�E|���n�����q�}d�iLi`���T�G��w#
f�cp�:�Wh7p�KA��YU�G��CӂN��Z��0����n���[��R��ʘf�Д�%05W�3G�n�K�W>:~�-?}�9y�&�8�Td�����N�<8R����79��L��{>�2��������7ܡ��V�sU��|�K��`��Hw�q�sK%j��$[���8q���0��*3H<@� ���a��5u�����o�!%@�5�l����7���G�S�gF�Ɛ[��o����-���K�"۴c���ܙ"�Y��O夂�bq��S����v	�UIc@(l�s�G�U=&|;l���"�<���2�`{��X��#�N�A�������Д���>��O�9�M�����eHT�'��ܙ[�=��d׀��5j��t/�Ѥ!,��I/�[���A�-хŢ��a����ɳO 	���Ą����7u��Q���sDk���w�|b�cr��r��AVF�oMr��(���b�+�Z
�8�3z��
���:�kTT�������>�� �Bш+>��T����
T|�7�N�qD:X��"[E_kh� ���Z�xuNc�M�>��_�[�&�(�1X(F��G	�ll��\ok��cE�N�y����������'�9i�ֿp)�{���yL#�	�B��6	��5�
��lh�yD;,{�����E��T�yq͸,�H`z�u;2F���
&z�8�)G�O]`�;Uy�gSz�2<4 /���_��X�(��C�h������6��,���{��*�B	ӟ��)�U��
�!6v`�����^I�1.<��=j�Y^V`+�m���~ǂ����E���26���L�u��ry]��s�2�(o"S��|�'�C ����Q�Z�S�ff��i�Vdu(���{����933���x�����>h�jz�7
UQ����8'��w���u��Ӛ5���-���8�Y�8Q�]\�Y�z�]�)���ݡ���\����YUؚ��I��k]�D������1�g���LR�Ւf� ���*xF����l=����Sz��H.�=�{�`�[mwK����4������w�����@��ӑ�g���q�d)Y��\6��n�5s�!`jf��$�$��aB��Tओ_(�O�|���)Z�h�@3� 2*=N�4Y�/�U�s��s�sKr��i+��2`�,�U'Y:F>�3�G0m��Rd����-`WW�'N)��Ī(��1:+�&�? �Ȏ�zH����g�Y�<��œ3�R**����>���N	~_���H2I�!+A
d@x��)��(��������w��%A� �$W����a%�R��,�[p%��~^3ߜ�犆�F�����]^Q�s�< ǁ��փ�ϡ�̛������2�m�)I'�0�B}�FW���r��/��4AZ1<VF����W�����r �������
�� �[�����#�"���\�d��`�׉8���ˢ���7=*Ú�L<��ݿ���_������weZ�;��lY�g�ɪ"d�k�T@/
 z���PpCY(.�)ׇ��Q[$B��@K�����۰Y"�~�4� �� �P)X*�I4�A��s���M�66NxR�M�b۲u�|�s_�������������Rj�vL������}�	�׾�5M����c�(�ad�M�)�F����k��0�;��e�Li✃��T�S)�Q��q �B�dX)�_�A֭����x{H)�
�����t=� �!�L�g,}xXn��Ӥu��Ͳv�zcA�ר1Æ]��JC�0]��4f�2)hdM���''Ɯ��S�|vKoft(�%��{VQ�N�a�B�	H��+��t<�W!�#emut�8β!��� �}S׎��n@V4_�5�偱��C�ޟ7ꒁ?�T���d:��40���U˥z�n4Ų'PpW.K�բD�����,��wV?@z��:��{�V8�M���7g�����;¡eM��VKT6� � �H�V���7dN�B��_޻K�7����dB��ŒfΚ����{!�Af
"-23\@��ܼ�L�Z1�@������QLEac`��oɹ x~(�c#88����9l
m�=(��0�����r��������m��J~���R��fr��+h�����Y�Q��c	�\�w��J�2�)��͒|�2�M���d6��I�������c����yB�R���{:���^dD�Y�4�$��Ç��_U|R�Gׂ~?�>_F`�-+uȿkF�Ӄ���
�]�����X6�H�x^�L�s �TrTthr�_��� ����F-,d�Pk��o,b�e��,�ԛ��	F�!����4d�u���b�v�Fº��Zw��:3���Y�3ڎ�SK0H���� ܲ��D����uV�u����MR���%ɐ�	�X#@n�i��ΕT���F�D�Z�D����G�!����I�x��L��/H�b�Mm$D}���A�"-3v�dm�SAW���Y��ק�VO�{���xxÞ�	 �;(�9�K�{��Ġ��~zp?_(�7Y?G;]klچ.�q |��w��DN?GV� G�c�������5k��_Ф�_2��nO�ɑ#G8��qӈ�o��ON�)ƢMN��吂sp$ ��r��)�x�B�mL&A�z�$�����a�C�*2��7oޒ?��?����de�ulb�U
t+����	�9X*b�)ݭ@�l@I�l��
�$�뻂_�I��ْ��dP�B`qy��UH,��@E�s6�>��g  <� gBAJ�bfy�w�w~�_�+�~�`DU �|�Kbl[	����'Y!?q�4���
j�d��t0	0�}��%y��o�#�>(C��l=�|�!U����TBL�"���E��hGn�=�3��VT|��ܙ�����&Z��9B�6ݛ�yao&uM"�G�����ʨ����=��wDTňK���,�^�fau��1���lOZ���,��_��/��qTtaC�5l@��kX�W=8���� w3��cTR!��ξq3%C�V��7Q]��p���u�:�t��y��� �8S;�����D�-�0z[nݚ��*�Y=$����z�{,��DcF	��lxp�B ����M�l��1SJ�Ç��B�D�8���B��	#֍A���7Vd��2#Bq	4�7c
�����b� 
��l�fK%��쟢�˱�z� �~�� G��s�����(�좦�fg?��O��`�ŗ���3�l�<�s�E\SJn�@ڊs��Xj�f5�DW��^�������%�s�8��Ѓ��ƻ�r.��'��)cF���S����䤩B ����́�^����R}�Bь&bʪc�N� �1D0
q�����&�@p(hQ18��C��3�$�D�p���scƻ� �1�+8�fY�&ӒП��K�n����� �V�����>V���:���xah�]�-������m�e���}�!E=!J�`e��E�uL�!��=��{ME�:L���Ֆ$����w�Z�������ɔ�Ú�����������ҥ���Ip���ʎo��8>
� }�e G]�� ��)�Y�O�]d��2A9<ӕ%�Ƅ�R	Q�����ڠ�ƒ�ݟ�S��↠��=8Q��A�ٱsLƈ����Y�����"��pp��Y�69���ު���k:�8wa�	c���ðSh�Z��v�y�-R�gxHm۶C^�̧9u�a<Y���/�vl������'�< _���ʷ��;�l(|ꩧ���'dvfF��{������^�����%�[����x�8�!�߲���x��Ɓ�)5T f&�&e��m
�Q83�j1�.�>�>�u
����پER�4���Ç��ѳܗ��+��g�>N�}p舂xU�S�c��>�	c��՝/��9�i���L���o���̫��g����ݿ���j�6ި�U�L-��lڰ^.]e��՞^��<ug�d�����s/� ۷o��nJ���\�8�8��9����x�/���F	њFU��'="�:�iH�F��M]���/�� "%*U�L�;SZ VX���H8�����	��J??�$`+��LDe����x6�^�n��{�؉m'N�S�<��B�*��pPU���n�)<�D���j�n�x�(K6ᅂ& 8�¡2�B{s�[��P'��8��6�q�@a�^��5ĎNR�J/,�q0���	�����n�0i2h������az)��c@B��U��,�&8�@�c�v��]����15.a�a����R��!���	�۠߁�6�kZ=pf�.�Y@@�B�20#����B�+ω��9�x�%ӡ�nN:!�Ĥǒ�7<���ԫfDZ��G��d�Lឣ����{�����"�QT�o��f"��h����_ r�ad�8u��J{u\0�q��4�np- @�g��e��~ �V� p�,��R��T���C�^Yuõ7,؍�|A\	Bw(��3�3k����iyϰ�)Ս�>0�K����
��ۊb�iFp�=ȗ�S2��; v�UY�h2*!qƺB�1gd��.�X�-3�=dK�Di�S<�0k�)��Ң<��s�<Ͷ�؍kҝ��w�^@n�&�Yp�R8��sáU�eܱ_}�;�V'�3�<�[��zz̎�Mk ��m���� ����<�ǴZWhy�[��hp=����O�����K�`g��ƔS)Ȉ�p@B�Ɏ��Q�]�ڬ��!���c4~��~P�!lTQ��'[�-���Χy8�-��L{�M�`�q[��>Aڛ�3�'~�T������9dT0�[h����;f�3@c� c��z�z��~��ȅs����W_�O�������8�Ε/��9�sI��cڎ{w���^Y`�WlU͵��N�����IJ03wg%�Mr�5¡	�<sx�PI��

������������k���?!�=��d��.���w	r�|l���/|��K��xCf�UC��6*�H�#���/7bh�LZc߼�Q#�0z���8?�����������w��{����I��fJP���+�ev��kt�$0�0%�6��79-�j��}H>ץ�p�(b�!c5Rpfw�͍= ��C�vkhI�A�k��:&���*!�7PM����H(�%��L.�M�����+��;1*�9�
�1*䨂#��P��h���D���m=��{�⍪��ȱ��=2�vN_��/R��� �²8��Ƽ ,W�x��(�2D��Fx�e��gC�qg�"C�Ń�@
A+�����a
�?R�(�-~�Lzp[���N14���	%y�,�!���e����X���nh�	Ѹn%���@?4ԯ���u�ˍmPi�>e�����mO�
fzF7P���<��<|5Y�Bd� B�~' �l�2����@	=I�f��|>8vJbz�2X�B���l#�(#`\p cD�Bk��b��T��N8֧ǵ�C��K����9�]{X[cC�ҋ���e��#�����*D���֡�"�֏��� �uEҒIv��9���"F�ܻ�V�7�jm3�hT��9���j���m��$L&cl<ӂt�U �w��g>7�	}@�j[��]��<*!A�C 
�����D6�H��Qe�F���تFh5�<JwC_�}IX[�.̨ H�s@�����uY��%����dı�(G��l
-��[��m�{���X�����m�P�	� ��'p��[:�������w��к��/I����=Q����:A������s>�1 �XK 	#��m5��b�W�.�K�:�l��	������0�X�a�r����5��$�֚R���B����	�����&KF!ʄf��׸�X 䚽��;1KhGNM��Q�㎝JwQB�DZ]���'&ni�� 7�@�Y�1�;1�S�틿������w�z�|���ٰ^�� �. �J��Ȫ�:�����_���g:f���i���Zg�Y�٬i��^}z�߷w���工�I^��<����D�]xߧ�yH��/ ���_�3g���B�T�A�>�1�Lg�X���9�=˧��Z֤�Kc#���S
���MJ㭃��SOˁg�����cG����hwݿ�\=h0Q�\c,�h� ��<����͕Y��Ӧrp�B�0}�ȧ�	���5�'&� b�K�^w�I/�m bX��B��<�g����ھ1�����L���D�I2�Z���'b�L��hT��-�%��<B�X���������;x�Zxa�6�!���{Tt�۶l\���וe�5x,.��C��W��EeD���%��yS0ղ�h�D��wHO7ʒ�J	}i�m���Ҵ�I�)�1ٰ~�̹CLK\}9��A�Fg�r���
���>Fu�E�X���xЎfTՕE�W����߻�����/�����H���kF?C��(6v͐���
�~��EG�lF7c`�ϑe��5P�L 	MDi���VT2�^�b�R*,��3č�Ԃ)��e��rL����cA(������[9�g?Ş�Hu�[�3zN��we��;H�<�Q�D�biI6��gv��d�	tr:�ZC�a������@$�Z�}0̀���S�8/`�'iS�+�8�?��)4
�0���X�>w�t���̈U�c�tF��]{]���pX�YJT���&[qC_�T5�4׬@>�K�Y.�kD?#�
�J�%�%�L9
Z-_�q���@��k#��M?����O��Ɏ1ꈖX��,@��
���JE3�p!{^ຍkD����A;����9��h�y]o|^�z�V`ǲ;�t1L�WT��b�.�Y(.+p��G{L^}�U���|�;r���ߺ5���'?%���ʱ�'钌�e�Z��߱Y$\r��q�^v�r�� ��A�`{G��:Ic��d�2�����݈A�s%��+0K��u��[��89b�K�fݘ�e�*�m����8�6!^�����k8�OhI�'����0K2''U�3�{0���?�����#��ꅫ�s�y��geE�naqAz4�z��k���l޸ɪP�i��ళSD ;w��B���8>�f�I�)�+M����$U$�HXp�bt�v)��*ih-\�.�g����{���+_�
���>�ӧ��J����)�֫�G8�[�q�Pܬ��o�;l�����$���V�kƨ0x��o��� ��+�}Qyt��:}B�\<��t[��JW6Ƹ6.�B�zQ�)ߒ͔m�79=30���iL a���U��ƹ3�A0�oSy�6�0�����N]R��	�N4A`�m�J�� 4����۫^X��
!�B;�����6A6 �k�?���c�j$& ݁�/��Pi�ѳ����T����rqn�����{T�)޹}��b]~��8=D4�ett\Ν�&�F�R� ��l����2U�=�����+8���8�R�+� �6�p�|j���ݮʦ-[��}Rn��|��wP��QUZ�l��yƵbU ��#z�]�9�=0V�rs��Ꙩ��NǭM�	/�?��	�-�&�`���Z��lң�lPܑ7D���j������$�'@P�Y�S�h�j��er�w�����������|�x�81vr�&������Ĕ�V ���b�ߋg ���fZ��n
�o��Zr����Դ�wa$g��YE@P���cI�|�L���=AJ�� ��C/�ք�A��G"bK��n�/F�;C����ft������J�°S�6U �ߣ��<@��uc�ږ�ؑr��&�Ƌ�1�
A���'C�����0�U�%���E��l�`�~A�0������C%�Q����\�Z����+8'xbQ��D���].������K�g�AJ�i���Q�S��_�Z%mz��*ʩ:��,��@@lH: @迯`d�\ץ���r�EW�~�%�Eb���[��/���<��K �HwWF����=��7�\N�:%}�]�́�B��+��$( �w�8�k�e��c�E� U��F� �6��BFa�닸ˠl�@�1g�S*������$��a�F�F�'�SV+��/2��`t?�w��KS$���֋Y�8$ PP�/\z��gx�Wd��\�~�i��?�aA����}y��G���,�PU�s{Rf����r�`���W�*-�_a�a[hH���,7�|x�;�'
��� ���#3 -�{+�� �a;F��	��"NC4m����˯�;	2��������.�Ϝa�
�����3iV6Ŷ����J.+g����}�@�"��|.h2���2;�,OxB~l�ܿg�&r��y���CC@�v�-����'(�ֲ�F�'���ƥ������g�Ѕ�T�BxL� �i�wM��Yĺ�g�מI�����V�`�jlTS�%�	��O�j�0qkq��L�r�:��a�}�����Jmq�GL��
�����3�p���8��6��;xz��sn*�=��'@yAi���\Xh\Ϥ�Bid�ZٴaH&Ƨ�6W���G�h��tT��w�4�uZ �����vA\3��LRjeͤ�����棷��%��/�A߯��pN����)�I��C��sm�G�ȟ#�*�Fb^X^b���%%��t�p6��Q�չ8L��T+m�ζ�Rा���m�w:�H�ij���\{o�Ѻh�u��F�C3��k(d���2��@$��t1n����	ft��rlt�L"ޕ3���*�(�Op:��&��d5�zT�4��`ұ�J��r5���Iwu����6�qjm�|
���n8��"eG� �iA��8}��*b"FG m�m�.}f�e,�Te�2ݝ	/'4#�͈�c�j̚�TjLi�s��rX[�'{���Ȫ!|h�9���P4;���(���C!B��v������:|Y�q�^��?�o�� ��׮�gC/��7[��[1����$�����~���h�9$u���2٤<���r��%�R �`���$M'n�� ".Q=��-�!�Zi:8���&Ь��H��R���Af]T�� 3�-��is�9�k;7��+P�H��"�B�ι�w줧ɟ��D����%��/~C�J�9D�h��	�KA��Vh_ .841^��i��Q��5%4�/.���,(��ؘ�6Vۙ���? D`�[�1�]�0�?ߪ_�̭���&�sK:U;vO�����H)�Q�ϑ��M��:;�%���ܾIcDM��W�����ܵ��앃o�-�w���q���f��c�
$���A�Od�8�M��l��C�PZ����T>�������P 7V'N�	t�~C[��KK
n[����.p�G���s��#�::J��{���/�3��_�G9����h�9�bB�Q#-�D����mVr�:&��K�&q��霱7��5	�fk���+r����m�e��%�������(ˋ�<�����V-�TOO�{�޼������p�.-(��%H�8�x��JP��Vc_�e���1�����?�p95����C��Mx��G�e�c�=��	�@��sJ�lӐ$z\[�� �ව�IaQ;$�V|�Pm�\Z)R4�;�-%8�7����{����;�I��O]{��m��{�uoܓ5�]��{��"�fT�0?��fI�=9)[9���\���M�p��$���x��h.�z!z�;��M����!��ʚi�ȅ�g�X��g�|H������W^���)9��)I��߰m�<����ducQ����#2:zMr� ~�aZ3L�$�{���d�ָ��go��,납��=��͛(��0�I*@�����+�3ҝ�UvC��ުY������fz��IJ߷��l�8,�<��9����(jN�����tCoi��{�����иJ�<���F  ������a�$x<�,a��3a�%���(o��h[-�anF�8-�.�D���N���Al�'g�F���f�(R�o&�1BW�zQ@��K��f�(G@PտWp"���;�K�eoF�ö�z-$YrC�vj�hz��e�(�D_3Nn��,� ��c�d5���!`�9		�|Ǳ}}#A�H
N0�ؿ���Qu���@�Aq����=�vR��ܾ=�(<u��	�y�Ny�ר�R��pJ˘ʚ��du->�ƃϐ��[	���vm��9 ���!�3����"����+&e�Mj@R�E@��p?�����
��ƈr9#Rn��P��^f��ڞ5����z��������f�"���fdv�� 8q�����?������_���Ї�;S��x��z�a�;��[�:��� �c=b�ܟ�S��P�H�F����4i4k�� ffB�ɀ=�Y�m�1aSB8�����q����6I���n��CXe����i��بk�$M����D��~�mE�t*#���_��ߗ�ߔ'�|\z�����fT�ݟ<~L��{ߗm���^��7`�f��m���SA@����9���e�:?N�tk�oQ�ٹ>�X�u�b��2M�rݽ4�4��)pK�����s����{�%���W�k���K��e~_��҂����(�Iv���sV�����9�R�~.�+�4nz�����{��y��b/mZ�A�a���Z�AA�V�}�<fx g��dr�TQn诎� $�!S�J���l�X����,=7i��$(Z��J=��}��p�P�u#��� 0-��B�N$�~0B�6e@�\gl/9�c�*��_�����`���!�#^z����U��B��;�����'����R��N�����{�uoƓ�I��Qڍ��#��` 0���b93��X�|�whJ�$!���{�Xy8R�с�DCy�����	&�n޼#�6��g��(k�u��:*�m��G��O<(�K�^ODΜ8)�=�G^�̳�oҬnA�=|�g0�%Ks3K�F�ʋ/?�.� ��A^�;!��(��y����V��W?��y�mS����w�\���m��=��c�����V9,E���);�m�^��`Ю����*+�e�.G&���'E�s����]c�z(�^%*{�~�m�l�ޮ��ܼ�u���0��e���S(p,�\
�\ ��{z�b�|�,�.l��ځͺ��ꙵ�N �-��X	�w|��Z����!�C�j�c1�Fؠ
X-lC��
\S.�� TVbŉ<�����dQhu@)Ӷ��Ti�'&�q�z�%X%�9���0�� T��C�3N5bc 	�p�����j�& �l�
���V� kmT�@�Tp�� �o�Y?<$���\�z�DIȢ?�o�LM���O<�v�~�}���Z��_��T����� �Ti��� >K\ޗ~�5��_��,LMȅ�qY�5&N���֗�HF�_2h�굧b�Vh���J�Dp�`�3�?�f=K� i��<,(��gdQ��|B��k�8�ֻ��В��Y��"�a�r�<� ��[�%/��"�.�zlKسS=��i�d9�W'�mZS�@^��*��Xk�ADNZ�V8��2� Ϻ�sa�iYr:(l���j�߶�<-V��Nl�o<�:���/3]v&Ƭ�3@E,�g�W��D����NP�vsB��?��_�aQ��Ҍ~ʴt.�RP x��#?�m۶I\��/�%y|��ʺ��/}YΏ����8t�x�~.�kE�!LQ�ĳZU~ZފOD`[\��L��o4�(�ߍf�V����|J&�f�����<�����ʡ�?$H��'_d������[ԍ��#!*$�F�շ�Q'ɰ�;��^Y)�#�\�����B�$�o��E��g���~���Rl�bR
"l0(���$�� � H���`�P�2�l�1_��	� �g	>���.]�]��x&��:1.�f����D�>Uඨ=ԡLP���/1V!����!�=9(�O����<֍���B�r��+
; ��5M.i,�3��71��Hw*�횜-����9��wo��_|��?5��'@���u͕ݠ4k�f}�q�v�pbr�ꢱ)'[Z�� �
��q"6[�J4萷\Bé ;��b�8)[7������iq���|V*��\�zI�}'+�{�K2u{N^�'���hن�C��S�I]���ȵ�k$���W~Mv��.{w�'�Ν�DBS�������ޣ���B^y�"g��_IR���#�蹱�x����}��G�+G�O��~R3׺�ͷ��j�8�8 _҃�W^�K�NH.�L #s3�򣟾��l�.Sw�<;�Z�BD*`�A���f�{����ۯI>���8:�	��pTzh�R۶�"�(�IR_���e�?��3VТ����
ök2h��ǔ�19��M�r�x]�I"/�Z�Tt��� us��톸��-� �Lp8��lJ�1s�l�if��x&  P@l�K�X��<H�c��o�`��j��ۥ�K�=� T�1�t:$�6����f�п�=�h6ZRH|p��
�0�O�44f\T�+r�ͷ��4��T@��26~S~�F]����ʕ+�VT�P��9.k��ӪH�ʃT�b���K�Y���f�=Y�7��|uQ�ʂ��Px
�uY�dc�A�����`��`ft��hOp� �=Nð��ŊB��4�HP{pٳs����\�ySJ���e)�e9q��<��W䡇��9�|{fF���ߔO�3�f�CZ?e��WIT��l��I�>��2㕚ѡ�J"T�+$t�8	���1�
����*"1A�j>Ȋ��ٖ��i"R6��x[�r���=�u�B�
,�~ku��F!9XQ�Oh��jf�c� 	��G��T�A�Fo��?��Gfd�"�\nʷ��r��9�p��y�����w�?�(��&}�=$(/,�4�	HB�8z���I���bl�����ѩ]A�oML]�N8��Ձ���F{��cԴ?#Q�у熄&����Ǵ5x��O3N��w�zSn��}�/�\~�/�^��r���o��?yB�Ks�̴J��iq����jW�@��c�w�Z-ۮF���ժ�EQ���� n��ޖ�H@���ɓ'٦��rOt����y��B�LHk@�mWX0�W�V
�}l�c�(��2���z9�z	}]�Jѝ��
�aB+G�n�ab�����<�Gh�>X��,���6�)+,/��� �_�`2C9'�ٖ'��i��..��<;���:+�������JZϽ�������ٱ���,�������?qc��4��0�=*��
)� W�Q���͛��Wo\��˜�A�R�Q���m����_�44��UR	�>E�Id��R^��k�ta��X��	�9#�ZQr��-�/H�tz"LNLS*�{{vo��|Jn\���n��}��q�z`�b�@����և=�9y䈜;u�����Ey��K~�������r�H�ā�����Y�0;q��<����{"�޷g��e=,���sϲ�v�:]?��~_/[U3�j�=s^&��K,��I[-�B4pȡ2��CFХ({ �+w�޴0b��<��n@���
f� �G�eu3Ԫz��6Kl���!cŦ��{m�`�N3I4rd &�0l��.��p8�G}	>c�LP��dB HF��x�2�c�]���3���iY�#�@������Bfmꁠ�̌�Z[֎P��.��
��<����S�'��V0��i+��:'��6�AC�M���=޶%����/d� 0�b�L3�G��z�)��v�m3d���)j&bw]��`A������A4!s���d��NP�lx���$���bj^3�j*k�kєs��ʱ�6H_F=l�1G�i������	���I0��������E�t
�È�M���^`%ah�N��s�N���8�>�<����ʒ��goP�5��]�� t^�%���_�A���kD��m�!ur�rY����cH���}�;�Y�Ќeӭ�*�~�hm+bΞgE�йKgr��c��UY[�!��-�����_�ׄ} ��=�L�����\�v �4�g�s$�|� �r�֎P�`a����9��=/\�b�g@�QYFo�Q�J���E9s��@�� ���Hg�8�m�����a�S��-ډ�m��ُ��TŖ���	p�=�>]<�|�|�*��ha���,j��R\�a' �ѣ�e��$�5M��!���� l�!V�P�E��ꩴ�V�:��
�	G13
�) r�X��U5��?��+l9�c=��[/��l߾�j�b�Oc?�\��Srg^��̜$�q�|.��p.��K�.�� ������$��K�{@���/�)3ى��$Έ1rL���9���撒J.�
�ja|��?&Fl��#��QﭢZ����	��QJ��X� =T�==��v6�&[��x�11@[*�H�=?�p����J��^��X�����m�S�'����,�Wo�eՃ��'�vo�����	��P�:�J:�b�%-��?^�M�5�p�� E��O��r��U��=�F�Fdb� 7Ǯ���g��ͫz0׌<��FNJ���_>׍5.;v쐍�3��(&G����G��� ��B2�e@�ҫ�PF�>	Q>C	wzf����~�i���Cμ?��~fA�t���ٹ
	!�F/�Y� ,��5N��f)��bd~����^HȞf&��g��a�S#p�F	Cx�
�/�g�}� �kc�i�=K��� ��KE^Z%X�������>J����a @�ԉ��L���)E�h])$�v\�9��&�)U�[�U�. x6��8�8�qN
���qj�������65P|31 �b|�('�"Rw��Yʴt�ֵ��5=[L��[l�TA�:a�S���������	���)�K�S�^��b�8Y�����F��2�Z��ݹz,�� uԞ���׮��� Huc<��l�M�5 ��;{�U��K�͟x��Gf���m��y�/�n�@1�q����1u;=m�<���s �zQ���N0�1�e$N�R���kz��ڍ������L��qڭ��[B3
��ӝ�ʉ���06�r����J�1ǐ�)T��}�+�留���v@F���_�}�UE�@,��8�s�(5�D�Զ��g�_�����L�2�����m3��Z^A�T]+҅�[o�M����j�LE�A�/
zX�Y�D���\K�+
֣�Ԩ-�L�2���Y��8+4�<Q�O\/h�`���U���i���[�E�ҏkFi#Ʃ��^�U�N������I@�`7� �0�v���by�. ��6�aӶ颦��Y�$��*��wVl��w�ն�ʳUZ�3v�C߰i�|���e\��?�3��o�.<�W�_8kb������@�^�
L�t&�w@DŌ(ڈ-����pr��DY��}���0�+/%~,'n�Y������Q�3b�6�r�1�Y������#�F��:�f�(��|<��:�U����y$�Ac��B�>����*�g����1A�� ϵEu��ZO�x�{�|i����^L����MT�ؐ���[�'@E�Eo�p_�3�n�:B7�������{)�]�ɉ$��p�g�MIA�1B�Rp����b�mt�Bn�������k8	��ӏ���:��_|��/z�˚��iA�#���>P4<.S�g���@�nE�ЎBb�����%��A��e��|Y]\?%44��E��h �ykB~���I6��k�#���3�xX��� �g��Tl�|��=YSz#B�����
vL�2sώQRiT�v�kR�$`�A�!�T[aO-�5�p��^n�(�
��V�9B�1:Cr1�	��qj[A���K |�x腶�퓳�1_
 zF��C�c&�������1��x$�yR���1���NhH~�[o-�{�G�d�H�
8��us׌��c_�	��P�%j�Ҩ�)[�}zN����W����z��Qp�!)S;E��@Z��"���1�^s���Qǉ0�]v,�A[���o���u��/���S�~�djX�c�����H�k}e��'�s�Q�
&�3fSq�Ѭ=�^>ZF�[�?>���wN.��ީV x:1��^OD>}�BݗB�~�6��3ũ��BM�f��.�ףp��ay��g�!"�)]]��:��_����M��;o����B9?d��>� �j5�*�f-�K�)ft&x:#�?�~�c�3��W��&�,q;��Ҧw��]o���.	��L��hg�#��W�ꐘ�~�R� T���lm��b	��Ga�Żb�2��!ɁX$�S�� ��${�b��=��)Xl�Qյì `H.ĺ�u�D�D�k�R�2�y�*W��K��9�E�7��Y����w^��*�Jf�1C3a����$�{`ƣ�3��!A	[)8�##�3h�� p�F��~����ye��0���w��ϴl@�1n�&������񳟲J���k�.�=�Ӑ��?�e���+ׯ���%o/�e��*���۸n�~�&�x���P�˂��H2��iE�6�9�$C,�q���E_� f��X{`����j�!Z.�� ձ�1#侷ʳjr�-��Y�{YbTBƈ~E�KE��x��������уj6L\�b;^"M�0Mt����/�,��������<�Nn=��sgh�'}��ҥ���p�㦻(����{�fK��<pe���Ps���
�@@ ER�%��m��n����m�z�K��~S�C�V�ՒLj"DP	��<P���;���Sf����w�Sh�M*A���;���s�5~������S��Rj~�$�����F��IX�qeˈ	|��E�N��	=腱��\+k�r��MN�����/?Md��#�4��D�b������4pIerzF���K���)7�Vɕ��b$k��aߪ�1�A�c9z�=zL������g�~D��B (�뮻���kؕ�W���syu����v�Mل6���MO�i����d�#R�H2����3Fk,�F������w�ec}�a�2
�m����Jl�m���Qt;.�<�\R�%fgd���ܸy��evnJV��h��ub}XJ�\:���9��&}G�
�|6z��D~��4v��И����ҙ��r�`�3>1%'N���(�D�i�:�[�q�)a69�[���"dB@�������^5�`l��y}_��i����1>;�J�$��/�Ct�&R3�8�=�gN�Q��i� �*�	Ѿ\Z�)��G��aj��'u/�B�������!�۷@�[ߕ��)�vvk{�>�JV
W�!O�X;dokSn��$���{����Y���?����
aV���_0��Iێi�ᬆ�S�� ��dUpT�ԝZS^z�EɿuF>����NP%����zFNk��7��	Z/�8^�rY����W�*����3���3���[�;��M�������lH���)��,�Hu;FbV(ET(K��$��X���.�P�ae'1��h��;d�E*��9پ���hMh�E�?i�[cc�7���*#u�����`��w�R�m^ +�o��/Q��``+ ���&*����:p����b|`7Y��U��Vu�+t���"����l�	<��iߨ� t��4���/!P$�QȘ�$�l���B���>F+^��ɫA:P�g={�=��X�Z`Ţk;�r9�/��H p� !�?����%�Y�u�����|�o��kz�C�]t�����G>+O}�I�9��P
ȝv K�z�����+���1 $L�r-X�*��18���$9��bz�ݍL��#v�U�r��G槵�>�@P&A��N�&1��M(Y�J]'�b�2dUg�W�:bжԁ�ʏI
89�0M�Lt���k����T�@�R�ꯝ�����V��29ч��uШ�;~;���P�fNf�(-�

������ʹL���2,v��z�f���~�i}p�U��Ǐ��LY._[�_׃Y�յm9x��<���t��!/_����@������2��С�r��;��_�7~����4T���!�V�l��{���y�m��ޔ�7��_Q����qC�����O�1y��3��ek�!����ȿ�W�#��w�gy�ey}]�����):�o}�/���#�ɣ�g:;	�>6A8�#�!����(�m=�]��n-'�Z�	��X��e��d�\��<�j�,_|������-���,5�������;dQ`���}�g�&L�=�6JɄ$�Āu�J9��!�vl�u���9�O~��2Mco�c�m_�s�{����O^�����$�B���/����E�׀=D4�g��T�����
<e���!V���Aʼ8�_��ْ�%�8!yV"V�/�#�9������[k�3�x&��⤩�B�����������ڣ҇�zP���z�"I⚚�����x^rN41t"s�f�;�{d]WZy�.����T)��k5eog����#t DkK���+n�^볿�R�r4J�8��p.����@����ߴL��g/Q��ĩ{�{(om��e�Dk�26�j �p�@&��Þk
��YZ�SϘ�C��KG���n�Lp�6V�GXu���G��s��UzM�c8���	�B�ӭ�!?"�$�-_�6Xԁ�'V!�{��5�X��ɉr��VԖu��%8l��+���RW[D]&���{� <޳׉=(�!���Z�, ع-늌�8����|ś�UȖ ��MQZ<�,�[��te�LJ���̅����b�,�1���}�s�̋r����K�U���s��2XM@ i�K�&J=�
��	�'�6,/�0�c@����D{gKV������_��%y��7�����O<�E�1�dswG��6���0�{��o�$�\(���I`O�f��(�#�������31ì*�N�Ϯ�8H�����B���W��.�Ī�(�2��qF�kȶ����8Px�r5.�f[�ƻ�wI5!.'�`�U�:i�[�Y8>9��a{�G���S�{q�|*�
�p�P��������f�H��1���O���l��b��MU���E�&z�ȅ;�0�(�ȥ��r�]G�/�#���\����}���4k9s��<�Č��o<-��"ok���G�_���dymK�@���<o Fo�I��(��ѽ��}��+���n�Q��W�1�D����
U*�拡,,@V�8��?�X�=sN��Z��D^�}��?��=�?"_�7͈�y��5Y��It�����r�����|�u���2����!#p_*�fX5�IW�:8Q�b��==�N@
e���f��}�QV0ƌ��������3�i�� #��xm�^�m`�l���KU��S��N��������tJ�%2<d�>8�GCA4�i^:t��gd?�l�}�)�&���=uzz��Mr��q6#>�� �  F�b�2z=cH��n9�5C�x���Y��c��'��1=�U۵S��Ih�bW:7~}�@�јqOb�����}��ɝ��;o���17pN���~s�F�ܹ��oW���R)�4�Y�{�����s���F����'k[�2�P��42Y`� ������Y"7M�వ�zF �e�}m�yH��{:�:�8};٪�e���ʚ�}R�ͺn,�K�h��g�g������P���ڧm�8�E��>��b���ٔ�W��[1ABiQ�·�l��w��S#
'
�q�8�LTP�*@����MG����	zL�f�Uz�58��8,H��c��\��S7Ϡ�ps����'
Ё N�������?u�eޘL��lg���wtD�����,�c������r'˲�Sߥ3d�dAJ�OE��l8^O7��$�Df`�\9�@��*-�CP��ۦ\B������?��^�&��6��d��d��bTY�_NH�`�r�=�N{�y���\�"���׮����/�\�^�B��$Ο���?m���0I�ƅ���OUOZ$`��t[� cӳ.����ت�X��M�Ξ��HXU�C�4�ǡ�����5l��w�8|��✠]�ό���V����s+cc<g�z���Rň����H�@�
��U�4c��k�@EA�G[���b^�bE?{���GR���+��������˟J���Z���ʹ�˃:h���"��`�z�,�l��5wޱ�9�tm��ZYql4��hp=N �oh�Yot䅗���<�Ȅ�u�c�	��YL�G���f�*����{'}^_ڒ��^���]R������ɘ�ʥ�l���]�W_{��l(Knh&z��u;��|�>�=5�?|�u�W�+Af�{���cSꠊ�~��XЌ� ,�ۻl��dY��?�˿� ��@�#�a��&��� nlr1d�E�z�aV��2������$@
���tY���~ڟ�����ŋ����,�Q�x��%���Y��򪝾����dGx��M_�g ����a�� ;���\�������?�^g�V'�̷��� �ns�*�.]���w�sj��q�(Ǿ?�2�y�Ӌ���MO�Q�osu��r/�eby0dE%�h����A�@��L9�
�h�Lv��"� N��{lm]>���F����:�y������Ƭ.Θ�?q�-�	��L�W���5
�
2�+m94[��H�ժ��0����=Q�@��d���g)�����䒁R����"�ȅ�ɖ"�^(����l�e[�ś���I���f��R���U�'�'�|R��v	$g�U� c��6�s7�3K6�H�%�V�^�`��X���
E��`j<'A���&����V�[���k�6u
�~�'0J�!r�bX���1/�~/v�q��� ϕ��oR�3T�����l����Aܧ���J�*Y�DO?A����~�,0� ������ ���;KZ���>`�4�@�F�m<��� �8:G,��c%J�<�4q@�vqI��# -�l�'ɘ~�9i���I��6UE* 7���D:Z��n�)h�w
�z�F����#�?��y�	VRf���\ު�ɵ�eR���/<�6�j�	�i�a�K��D�ɥB�=���b�"�N���t�nO$��x6t`,�p�v#�^�Cl�&!�*�|.�ek|8�&b�6$�U�K�Z.HP��R�#�eu&
:��}�Ɂ�y]����M����݋{�@"��$S{��U��L�c��j?�^U�������^y�_s�u���ј��j�$����- ON��QWS��FU�Lh�p���29����'ٓ�u�krrZ7֞�i B�{y��Tcd (kX��GU7v[r�Ɗlml�h[���<zP���\^���@�t@�'5��ʓ,/���^}�@SS
�V���9d��)R,��}��Eֶ����Ĵ�4��[@~W:�k�eC(���.s��b�6v�l�=���g{���b_<�)���v�@q9*~3�)kD�����)��'I��ȁ[S7O�b�������gx�Hu��"�`B�P�a�'0lB�N�,H��G�D�!��R~ �Zp�b�7͢]ͪcW��j����b�Rld����&I��(}����u��4�^�SJ%�0�i���w���u��ٷ�;��E�������r� g� ��� �.������mZ{�\�������䖕�� }�T�ZRs�O�r�޾�yҤC����Id��p��+i ���9ɛ�f�V��hK@����y�fچ�)Grcm[�.�gZ�:5}�#lnˎ��50b�\�F�S����t	E�@I��^��=[MYܬ�͍�,o�L��-��,�m�ْ�?����On?q�CЧ��c~���}Ȫ*p�e=SSS��O���MV������#�8�q6�����q�4�'���c��v��j)b�lę����)|�� �X�����>�ؒ���b:u�6L'�(hI�׵�:ub��T��zm����* �0����9�h�P�F^]�f��bmx��K�F��
�s<{��5pUq|�3���kĵ���3ND����Iy	p�왲%��X_'��F�7��c���kl&j���b�l�@Jm%�9z�οX���䣏>"}?*��R�q�v2l-CQ����]�����ի�����̻�l�1p�8�(��Q�Մ���u���h��<��H+�w"ת�}�*! ���0ڎ�I|���f��
  �ܦ���tQv���\ǲ��*�˺O�Z�t��)�z�M�J���o�R�ى'u��T�.*s]�*���4�g��u*�[٨��vm;M�j��S�����7�������_��i�~�(,B
A^z�z�y:�?���L[C���0+�8SL��[����E�*��s�2�A��xd�������x����)h��-���nׄ栍Ӷ��$�ʚAK�T�N�d-�D�Ʀ�<��@e��w������0]�1M��#�H�b�^8�0���P@�oU���1L5��h}$.�]���%Tbg(<��_-�KE��ڀA���B5s� ��	�n�&�f���gw�df���l��D��N���4f���AG���0����5X��������U�Ȓ�~/"�^������4 �5�����4$0z2�*���%�	@4��tɕt���A�K�Rk�A�	8����0</�ɩ)
8W��@�].�kP8� ��Rn�kcݩ�@��G@q�ᰥ�{���K�g>\V'�G��΍�́ B��T���g����\��b�%��ʸ�
���a��-mݗ�h*u�@^'e2c_�IL�?6��F�-�s�J�c�ʎ,�Vv���l��a5�K���jۓUQ�|��7�9��*�Z\#�52�z�AQ�iڄM�j�|6 �B%)116�M"�S7��E`�O���T�/���L��M�ЩD&Jɖ{:�Q~�v�AJj81��}%K���s��3H=��������8�l/F�0��������	R> d*Lg&��7��A�i6�|�*�'�!k%'L�xN0�骲���J��������X������m���9�< �\ �Խ�B8i�gSY�O%�
�� ��æ�>˓�m8l���N��ΰM��nJ��I������/������{��w�⅏	�G���o��������y������r��T�g4���/*5=M2�A[m��N|���V-4|
���3���5��jG"�V���q�$v�V�J�Bbϛk�a�PF���ޕjI��ڛ�F]"�}�/���΢4�������%�[E���"����y%�L  ��IDAT<rL&�J�4�6Z
S����7��.��pn��9UȐ����ږ�+;�O|�G?��7���|���YG�g�>�@��@��|��mR� �"�)�ݠԧ��)N�,aߕi7��A���v�FJ�Ca�JP���*S�UG�S��LA722PM�H��ؓB��s�����[}F�m}h��e���E9�AC�P�j�SA]�r&�)��՟�%k{Ү�W��=$�%���N��UC��������80����E�p߃H��9A7�GΰA���Pc��ς*��0���I]��]�H�^�%G�ׂ�ʞ8D.�����%S$2\�P���2d9F<���BwаqKz@�����ґ�y~�(��lcص�Q�����Ȍ!��hi�̭��	Q�Ʋ#����Mr��89�x����］�0~��5(�{��-�zTh��A����7V��A��R���G����+h����a!	�<�
 [K��nr���{�;;�����H�M���Q8�%��.�!'���%���Vm�T�9��m� �~ԕF�jΪ);��L�4x�5PI�T[��a�֏�������& @�w
j-5��l�5���Uަf� ��&gef~��ա.���y�3�dP���I��vs;���C#p���bs� ~�j�=�]���1`+�*�|��	2k#*X�p�{6���7���#آ�L5�
K� dS�L���S\�!Il"�R ��s}�d��4c��`ӄ+�D�h����0Υ�+G\�V[�h�z�Dp�8v�!���p��M�Q���)��7�>id&��H�`2�E�qc�M����8�r���t[8�#��Ȓ�'�bWÜ�k1�"&{��&`"(�D��W/ (ԑ���F$>��E1�v�1��)r\CXЀj�Z���eyuw�	*)8�h+{Х˗e������ӑ�&&e�\k�Hpvߍ�'�ND�F��|�����u��M�C&��!M�'t`q�/��4u��C�
cb	W�{�e�隖A� ��(J1�h vM�Ύ�<~Dz3���ʸ�ג��v�ؘE�vIN���M���&��Oȱ;�����X%��Ą�J�1�AC�!D%�-�$���m�������6ޘ�STP�Ô	8�D g�}}�|.P��XtBj�Ao�O<^%���q2!����18����=���X<t�;_*d쀑J�F�j������P��u���ó�9Ձ�P՜X�4�����26�@����p�A�4ؑp�=(���c���8pB(� �pm�_BMh��^-`���z)>��@,�,+C;�Z��ȱ�����������;r��1����}9u���J
��(��L
�1d�Va�9̈Fں���ʲ�@W�n:D�7p휬z&C"4_��#��؍��yY:%r5$��6�����/n���'>xp����v��q��E����Qu%�Q\�U���9B��=!�³甍���͏���3"WT�0z�`�	�2�|΍����Rw>����259N��+�.X���P�u2�,S�&m;'sL�4�{���'��0Ua��y:_��a��`,Vc�t�Z���nS����w����p��ͱ$�����]��{�+���83�⾢LǺ�����׋���
�v i��cMA���V��lY�DT���{��^��th��=dZ��@ڹ�}�Ъ���9@�: ��7�h="'�Ma`#F�'q�`/���S:܏t�b�j����K����D�_c�������"�����}%�Ԟ�*jk`3P�C����YmM��$'�GF��nCZ�om?���l��=��zʀ(2M&K�i7�h��M��Oև� G���0Csb)px��M����=�k�@�/�U߂��d\�Q�8�DLh�m��*D�*H��ߏAgxs��lϢ���<v/��ԁF�@ϼIZ��������P �LnSRPG{��e�Aa;.�u� +�h��:T�UP%�*9r)4�g5^�\����F&�c{��5L��%���MÑ`��vF���h2��(��2]>(����|�Ow����j�ʲ��$L� [U���lۉlݼ�KԑC'Nɑ�����Q^��%ظ显"�.�4�J����}�V����ܡ���q3���,;�e0z�)({m��;���G����{�XƧ�X ST�:3��&��c�nn��6�"p����X}?�;�Q�S�?�_�^�u�� @�-�a�;\L�`*��'�B�fj�.�T����Hi�C�\��bx
�@U�8�Nׄ����Ǩ�a}8u�Z��8�^N�8N�9�C��a*��Y.�x�W5�͹q��"VYx�~20��ȩ{�g~�K�@���{���kW�i� Fڵ	���*���^&�[w��\�g#�����Oj㓸�ԦgRf�	��u�L,�N9� ����ֵ��*�*6a��or|J�:u�TP)��>��-@���sE��C�'�P]�v�l����<��Jv�(�Ԍ�����\�rT4rL��jPȱ���������]��Wb��J�ǋ����K����)B�>�\���	�%����Z��Ա�ƫe�>>���':`&�
�_�2�`�Uc�Y�XB�9)�R*C�<X��܃�n@;T^�^AU�HaWz)��͠5�h�w���>�j ��a�v���}�g�A(^ ak<Z��z�pPX[:�" ���a�}�5�'��B��Ra��@F��UK,04Z=�v�q�}o�U=PA0U�a���Ģ�V�0$��&�qƬ:�,�q��G�X5�D��L�#c�6��g��Ԡ�En8��q�CjK��no�I��Z�K�PK\H������X���9�����`U=�ݠM�R�?T�rĵ����*@@�*]V�0�z�{`�Њ/X5 ���I�OsĨ�hb���,��sň��b�ɑ&��l��|U6t��o �-��ֵ�ڑ�>����ϊ	1�j���o����ɜItDu z��#���i�[�;�3��+0c���h���H]�-�qT!�<8�ijvRܽ$2�����1�K4�>�%h�u6t�HޫcE�����˒jBrhaB6Ww�ڥ���#�?��*�y�9Y��e+lkg��sn�InI��6d|jF�m~W��e���:�:��m^jȺ�MIF������%�R'��.��{q1�r������O%P&�r���A�4��Vc�*l��L6�LC��.��)GQ	��SL���{Tfl�z�&�)�k�%G����SO<)?x�U���Y�/�s(��z�"GvO�j�=�ޢ�u�����H��3�W/2�0'bC����/\��M]�x8���'zԢ��d��kEn?qD����5�< �By`O85�ȎIU�O�b��y�ZA1c�F�+�R�ݓ��<�%�*8�'�7��a6��
� ��A"�0�9��+0�0n
��%`�Sܘ�+/ 7OMNK�Yg	�E�Pb�j��9eӢ�d���jm�5�sq.�a�����4�H�H/�T1�5�;z�p��=�ұ'C�'�4Ba�`!W(d�L�`0��	(���uf�0��~Pfg�X%����G�/Ƙ�M�檱�^?6Μ�XΞ�Pv�73��ɯØ3t�}��VU �U(��g%�vG���	X#������`������=�VӮ�Þ��Ĝ	��[�M��P�n�o�2@�C��&N �@�,ͺ�r��D7�Y�UV����V�((��efb�lb�1f�o������Q$1�&�,g�̵�p�`wE�@�&B�DdJ�}��P
��J›���L�U���`���O�Gw$2��H;;��Z����K��(��̬��5mRX�G�X%8���&j�=# t�~���9rIa.���^�˜�x 'Np��܁]S��Kˈҹ�@�G�RHk��0�$o���q��֚X%C_Ũ��� a�1[�}�j��D�ڍL�n�pW7s?�nϻ=	-7��啌84�6ehjp�}L�m��U���bɆWE�^nB��ߓ|u��g4=ke�KL��p��t���{0t!�c�ھh��2�e{ͷ�����r�"
'yb1=@�.�S�vy	 ��/��V�jUU�O�RuevzAZ{����$'M�T� {kM���� ����HN�yB&&�����r��e������}�8���p��������r��{�:�?� 8�T�A��Uvp&A�Z#��Q����jB��/P|*���#���q9q�Dc9�����w���,
@Z �8��g�$z?F��WWB׻�ݵDR�]lJ�r&\�;�����c�|47�Ӣ�P$�Ɋ:�<���t���ןC9Ώ�b��$������7V)d�A�F(En@6>�U�t�5 *��Z�
�� `ʋzX�-����o~�#�������`H��VO�-�и<�j���e�Mwx�o��Q�A�Go�X�r�\���&� G>��;�4��
��(��~��g?;�A���toc���I��A �!��� �]%�U�0rU�!h6�T��:K�)���A����~fj�ZB�r6��Ǩ��D�B'�g���f�<Bfj�m�O��M�t�Jce:���/����;�fFE����:�r�z�k	�0-�U��ޮl�k yU��u�������4M�:e;q�\���^&���dZ
�\�Z{�R��^�d��r1~Zo
�{��պ	�����^)X3����Ѭ[B����d0<hS0H��(U�L�[6���$�8�Z0C�6O!�K-sD�f-b0wL��[��MA"��:"��Ȃ�]T�d_3��+5�f�0$���!�%V 5
���%{o
&�"f+v]Vݱ��?�ud���6�xHļ.$��W1K(���$·:�"+Gi�j̌�w4h���DIձ�;�;���
�!L�����C��A(�1�'�8���	ۖ�������u� �����Ջ��QܽV�B�3�9���5�")K�g]{��7���
<���N����z(���E2�;P�&�+�p���TLz�ۢ7��Չ��!�����*,Lb�MSN��	���(U2{��z��2F��? �5��`FXJ��b[/�L"��+�Jq�CRBs��5�lj
�9I����5��ξ��l���¤&���ձ
I�v5��_�D����c��;NT���r�;�<>%����\�.��|u����rM*S�5ٚf"Xo�ĕnY�Vǡ�-�6w,
�B��Kz�>�(-�{�ϧ���*H'�*������}�`� I�l���f�4����T��3'�{�OH�r!6$���)�6.��M�I ��C5��%5r�PlJ��+�P@�G(mv�pQZ,J�\�8"g��"���4o�o���b)����r/���p�%r�DI����؇T{'ǋ��:�d�K�阥k~f>��8���+ʑ�ez�Bv[h֏k����k��Nrs�p���j�3J��)�t� .�e��>%�f�����q��=��X�L��b?p��4w�ׁ��t��a�7}��e�B�vh�ì����||��/&�,�iq�ę�7���*�d�8�5�p�+�(mq$�@���赎M�y�}���s�]f�[P��Ϸ�C�*nI�4���������n*��}/��W�⹳���ѣM�M=��zn~F�F��jd �~賝��eS�uO�����%�V]�_�J��12h�iS�Q��X��kb��WV�`@��A���:P�i�V��_���i��1�Fn
�~�	d9�,�� L�5ɦ�2��칧j\� ��u�/1���i �{�4[t�e���_���u����g�N��ݷq^p!�N�huI��v<n*��u8���q�ڊ���e�	3nTäOg�"y!Kj@�\q��@H��@:`�P1Ep	hr��UNs����*'��9:n���v�g!MPoX��`R7����a.o�)�v�9u�%TȬ��d�}\5�X�0c9q�L"�L��,c�Ɋ�:�1�:r���Q�Ѝy#��m�Vz�N�v��k��ϕ�X��˦�0�@@3����q��|o'b��I���3�C��t�p���b�Z8L�в/�Hz߃�+e�h���@6*z�=���/�ړ��ͪ)�ѵS�I��Y�
#���[��=��3
E�m�x9��B�n
L�
~��OR�\�瞋\�0_����{�b��w�71BMh����v��l�ސ
1:r`�Q�G��x�d��>|�6�����˾JE�|�!5{���LO��&婧�Ȥ���[ryq��wk�df�r۾��w��64���a�0�+=?DP���n���N��Wp�~y�
���#�@5�ZuV�t�O���P�s�X��2H�b9����.k7����y��,��m,����{�]���ԯ��J#d�jo�l)�]����;O�'uQo;�Yf_n\Y�K��dys� ?��&�ԙ&��Lybr\z�q��ܔ�w�.Ǐ���?xY��GN�8�Y{8�����2�̺����<��G��{�ep��+W��w��w���A���C��3r��!����������}O�;��ۼ<�ȃrJ3�㷟`6 ͓����@Wl�;���k|X�߼��{��I���W���}���ؒd���֙*'��3
�"Ya����F?�Q�Բ/���$�i�;��1�
 ��8N\�Ĝ�� ,�H]�^�.���`���gF��MH뉭|�-u�ŗ�
���F�f	FfѢ��ە�٣�t ����Lݤ�d����������`A1��yM�x"�$�;p��������t�Ξ���q9�����c2�Nybb��$]��"k/hV�	�y5.'4���������>p�p�c�6���9V-��Ų�{{�� t�u�℁���I&����<`D`���9��ԈC����P�W���4Aɜ�8�`�*`/����b>e/��Z<�����KfQd� ��l���2��S4´��g����S�ǦF��V�#�MP���:���yS�F5	�/R�9��:W�!Srd�KnD9G���ib��Sώj�+�/�$�S�Hl�x���Km?��&�U�"s���M���k<?�Ǻ?+�D��15h���FE�W�d�"_�d�+6$���9Bt� ڠ5��rna�<"L�& �(C������4�h�dg�qrh���`�!8�N�*��F�ka#�!G�}EL�	q�1�>����=hQ�Q��^�A�����4��lg�f����e+a�ө�=�g�g1!��L`m:��$�C�:����$�qa�:��`�6�,[�ʤ��@��Ń��	p������g9����j) �Lllrձj^��~Cv7�dks��ւS��O=��;&�kK�dx�qh��b�6e}���L����k;[k�#
R�LI����$�;29��-�Zrq�J���2�~���ҋ213'_��o�k��%{�h,�lH!��]V��vLn;�_v���5ڬ<N�b� �R��u��ր)T��K�~��㑁��ק���en�I��ҵA�Ֆ��9-�c25��c��F�s��)Bb���q2r��B8W��2�~?n7������<���r�2>&R�i������l.��q VΩ�<��S��F�ё	�l��Q�0!;o��f�K#
��n>��͛Tc�~�+���c�N�7~�K����t78�3V��� ���|t�C��{T~����s�g��W����i��?�i��ܠA�l�Km{����Ԕ<��cd@���ՠ�:pX��W�"�Ӳ��A-�	�L����Ԩة����:���?/z���d�U�U���ٌ�/~eyLP���}�{�Qk�@�Ĭ�*,�?y?682)�#؈�h��W92b)�l�~��=~���-S2���.,w&�L~`c��)@�����ƺ� dwMfU���H0������ ��k��nC��3⺹�9�ʯ|�SfV�WV	��77#��=�_�9u'��9i�Tj�K ����!����^��3��SF�?7/�xFv����I�?7V0��S��{���}t�̲|���6�Ɋ8q�|0i�YF��^�����g�|�ir�rѲb�H�o"���T ۓ��Ā��8��C���uh��3�xT0���ε����K�j �5��~:���C����D͵�Hy7~�  {���Hrl�r!��T���9W�^��o��Eq_��&��w"s��T��?�oY����9��<p�Vݰ�9,����X^�ǥ�vj����#����[��z!�ʝQ#F�{>����5���������t��0c���	9���*��d}�1?�I�8��+V6g�ݐ���:UV�����#�ۿ��LҰ?���ꫯʋ/�h��jaw�m�i�h�6>���r� �*��>+vx�Է���L�R�!� �ɉ��D�;�8�"�vj�k�Y�9з�A���~ ��ePHE��NQ�\�V��)�W����Ui����/hP�!��r��;eF}��?$��F�%T5���u`>ս0=���������W�3=������&��Μ��������|����5{��weߡ��,)��$U2Mț;������2]4����༡bi����5fJ�|����T���(\�r9����1Z��>�����u]�=�h CB'$rj��IBc?�S+Sb��8^�;���=![ۉ<�Wߗ���:��SO��?w���?,�=��lo�����rmQ�4�����4�n�!�L��e?\���Oc;H�Y^�!���_���������></�?�����K�{ꩧ�������,7�w��/<�yY���<�Z<���>$O>�|��/�g�ǂ/|��~ƷYzj﮻O�ç����?�s���}���ο��^�rI���߲܋���ֶ���O�м�1�0�ZOL0�a����u�lðD�9 ����ur.]�0��^��P���!�SV�����+u-�Q�Q
rn�q��[Uf}�3*�6:����	:� �J� ���^g /de�Moe��^m�Jf��w���F�p2#��� �u�]4���m��{b�@�{�C������Aޗ�C�Y��"2]+/���O5&Hu�ЃB����w�����OL�6�n��$|r#��Ifl�� �>��}��I�������A6`P���)yH�!xg��74���kϟ��J��4�Āg���ˌ3���g�'���:��3"�O};�,�ЀA�X������]��A��K�$�	P
�����@pNb��A0j!�=�̔]�(��LRص^Oj�ئ6R�c���#��ƍ�n�&��K��U�%>$�K�R��[�Y�uNOO��{OJ.��b�,x���>�Z����x�%�\c�s�>"������l����
1x��_�IVh��]�+j�mMtD��[`��c2`h�%/�Ž���p\0��M�%'~�������������7� hP*`�oy�&eHv�6��w]��}��ɜ:���3�	�1���_���n�:��#�}	3%�l���i���0�^���B���V���B[��M�r��K4�ؐ�W���0ɫ��&���56V����er�L���V�c�n� ������%G�u�lB����r��QV��/�4PA�|Z��|���؎7�<�wk�g��w>�F+���u}�5NJ�g�KH�0P
=?�=o`{qC�����f�9^��6��ގ�X� �ʹ���S���J��2%�URWN���H��8"��璞�̪�?rd��W��� �m͠��졍��c�2�?w�
��ܕ�j�b��]QC|N��)n�@��oK/�9�2==)���r� ^0�P��
�{�~ +��s�9G�x�y=�8<?��O�~fy��h[�y�-ub�Rx��J�����"XƆ2;=#�>��\�pQʅ�,޸)?|�%����rH ,�Q�@�T� �b�	>�fowxhL�d�=6�@ �������@�"����kff4��ҁx���;�[�LܦB<�0^>��糟��Ԯ��
��떯����y�~(�v{-S��1��1.���n	������^����+(��>{���������g��~��%#|�!��i\��A�޷UY�� ����ߗtƩ��N9��Aq#�A����+{�Xc�k{x�Ԩ��g�����׏�F0l^�DJ��.o�U�w�* Y�~�3������4??����lq���)������>�-�!��Fv{�6'���@��=��긴*{��`t���}D2GE�VĄ�Ud0Id��<1AA��0®��I����M�8pb�i�YD]�D�ם`�U`��#�c�|О���\]�:(� X>q�l�� FX?��p���w{�3H|�
(����g��׮� A�)�/����f�42F�Bq�E��&���l���+�*$%DU���`�<��}���y��?��?a��s�ꏯl���)��Y��{U���Ԭ�mn�~�gv�E,b}b��c	�ǌ���mG���_�U`|��[Ҷ�k�L}�隰&d�[�'�˦y��􍓃`���@l�\{���4�N��L2q��bI��~�ӏQF�zt�9u)0ъ��/=M�<��uOVe,��O�F��͍-^���HW�����]â㔱)4[O�RN�U{����I�۹_~�'�:������˩�CQ������á|xaQꝖْ���J�2e?�LE�&�ļ��S:�<{�=�i����a��	�âh���+��*4�|^�~���qĖf�8D5���I��B��lPQ�F+�!t�BL�-�����tF������)=��� w�(���p�Ѕ�goml0��� ���UP�nv��h�,���d��7�Ӗ
cҍ���������@
�_(Xƈ�/��@�4�M8��N�=:0S4ƁM����Ѭ�hܸq�yvvޱ�V� ��@��S��a�ӽ�s�+�%�|2�����|����s��𯬺�p&R�k�}aR��NMu�	i��I._��s��g��������h�ܿ�H58F���p<��,ˑh���� �D,hC�'�)�S�` ��.XT	�5��g�<y�>�=��ސ"� �`�`��\`�^��b���$)z]�d�|�h�ژPӌY6[q��3a��0��ܑ0#(�(e��͐}v�\F�=3ۼ��Ո�Ǆ~��h�Z��e�v���hwq4��9|�{8���������t[�OS�ü;��f�^K������.&�~��e�Z9qc�*���x9a�S`�ͱ�r"F!���nz����Fl���ce`T�al��}p��Y�:�Ea{pzrJ�W���;G�ą�J�J�#dS}p��><KZ��ϟ#F�(p�H�j�u�U�6�1�k�u:��*�)��1�� ֦}E��H�J�pc�U�{��u�,���l�¥����������٨qS�=�v����� ���|��������b��/�a����h�X��#̒#���tI5�xb2~�"Pa����ձ!NYc�1q�S�}���.r����ae-6��L���[��R��&x�pM���aґ�srϩSr��Gr��������ÇdU��)�r��aj�C��=��-ȶ��Ѫ�)Y�n��:��@	��h��-Cא���{�����Q���Z?q�<�[��TU���,2��_&�겴�+��G��.���c�'0��?��G�e5mG�T.�a �:_.Jk�u L#���������,��cG���,ghW	�b4�!�_�!�0�@���d0���iuF�zO�,{��`TԹ�.4X�����z��'Hz� P��F_`�i��`�^�ղ�
\㎓G������`����t�<�-ݜ`>�1�ρ#��z����Q���V�����m��6�)(���ntx?�C6�`8q3J�Ǎ0�W��k���_޹���?+H�$M���?� �M<[���J�M��Q��F�=hӦ��`<T5����b�}Z�/����6�+�]H���+p"f0}f�fXc �:�/�Ev����ׄ�uFxOlg��ApW,ex�OYppxS;���9�Z�鶄��V�b0������� ��~����5J�&@K-N�A��!�VP.�d����g�p�h�A��O�@���+��!u��'����3�M�ὑ�1sO�̱�-���Y:2m���D�X�F�?��s"�}��/MS��El�!	!������
���m����L�
#d�2�|D	Y��iنH-iJ���?3y;�����dYʕ�#p���Ȧt��H�4v����?O[	}*��>k�����z\��F�٥�N�QK�m�Js�Q�﹏���v��c�E��!�܏N�yۀ�
��ױ��W�2zܯ�rN]��.��;��`��@l�ۆչĴ�����3<VUI�T�㉡Mt�"#�)&T�}2�ٜ��<��Ze�*8����,h 53�_6&�Dj���wpeR�m����[�_���gc��̰���Nԧ��?�����2"�`�P�21ݭ5�򛨎��3'�#�&p�-/�	r�^oY��6�b.����ΈM�Z'�F�~"�����ק�n,�,�9�3�p@N�AQ�'���,o�0-�
y"up��n�:O39X�*8��g2�dJ��qsyEN?xH��!"�(cS�AS�U�(pK�ȃ> �^&�Jh�j�e�^;a��N�㖝!���?�Q�f����'"X@�C|,���SQrK������t��F��r睧da�u���b���O��scq����x������0j��lN@�؇?�����VNЎ��O�����Il�l���k�`R��]LW�?	�|>E�K
+�bA��12X`�C��ӢJ5`.����ϔ���;��@d�5����h�3Z��YՎ�G���Z�GD�HyCj��b�X��~����Pj�"rp�X��7����:�Ё�Z0	�0?����������E�# �>]����� �~A�����<!���b��OXI���%��K8��ɜ�I�~��������u��É�=��wi���c{��-������N΍��gF�k���r㈫r��CcLUUnK����0��,����5ìt��>��i\�ic�h�F��:s3�r��������UY^^�u`T���q�u��D:p���i7���������ǵ�]g��v��F�mj������7��ח�6m��>J����a->K8o��$��&�S�s�Y�*0hKWJ,#s�p����g=�{�X
���:lI�9����fV�t�a`Y�s����*�A36���Wnm/E 5$QcD	�嫷xO%�v�Q`qv�t�L�3�/,:��р���t��ؔ�O�]�VM%h$��V��Iޜ�.�YE9 N�	pRX�4o����@(�/LW�A^��C!7����n���#'n���<F�C�Ȩ(��w�^�� YZ�AX Z��'��j�Ve���._�$�.\��(󲻽%��y;[�{�kvտ�~����������9BK_eO9x{�vk�KC�����K�z��+���Ծ����Ҫ:�L�a�s������Ma?	�¡��Gt4��$���F ��K���Yy�s�s��{M?z\�wDv� ԉ��wߗ��<��i�wOvv�Γ�����+/������ ���u����E���KcS�, �����b��n�{NN����g�\�!���i����r��u�����3���( K�5�@�e}sK��{�K_�ͭu���| '߹[����������OMj�sR�]� ���:G�@�S˫3�Z�<�9�6^�eơ�$�Sw8Y]�9�p`�D���Ӯq�FdN���xܐg�E`h��A֞�6v~"�p{�v�'�'����5����I|�>����`�1W̹�t׆�3s�擭��.0x0�xMLNp�����]k��8!;�,�~K��wx�@n1��n1<
�K��^m��J��P����LkƄJ���Gto�q�1�X@���_ϑ�G,�}�ȣ��̗��˕"���zR������|�\�z�e�3�e�Vul��m,��v�
�h�0�Ve�O��<&d�k�^q�0f�i�e�0����'���qI=X��P[�h�t|հ�<����o��o��<��_�������^o��D_�c��Z7����XRl�C|w�UTb������E�P{2tc���9��3���N�9rU��q�$���E)�j��1����ʍL'��@��Ks�u.5|�~�}���_��<��Tȫ�v�^�>	�,R�S[�+Z0I� ���Ȧ�a4�h�,@�hK(�6��)$&`��VU�v�c�|�k6��믅�襍�S��pǉ�x"P����o�s�='[;�,��A4,7�5@��DbZ"�4�j�_�r�M� ω=�����f�&AV����R�B�����N��>!�C� ����~��OL���{L���{������H�a���zm�}2qk2���T{H�{��V�d{c��*{}Y�~]﷢*O������ O?{anV�_�DY��2�kk�pf��kW�SN$�:Gl
�1��w.��!y��z[%%�o�>���.v؎��t��������A ��ԀS�hl�!��E��IX��������×42l7�������3���S��S	p^��fнXj;�k��*O�͛���|W>�ģ��G?G^�zS����"{���1�7����uz�|pv������Ы7qo���08I[]��Mu⅋7�21��7���Ǽ��O��ӟ}����4#��O_���9����.����噧���>����,I�V�ʍ��W������~�	"�:�����r��Mp�J[��o�/�[����.�0Pa�;}�a���ӅȚ��	8G\�%5�g����	Y��ΊZDn��L�2�F��j�(8u4��k��6��G��@F_��0� LLR ΐ-���� ��}���y��1�&^4��JP�p���9#��=]TU�9�\�v�����ӑw81�Жuw�r*�������϶֏`�$a`��O�w�"pY�\sAO��|T����F:}`��˯?���'� �8���k_�
����達nc}��v��E�z� ��W)J�/�~���=
��"e0�C���ܰb�{��MȀ��	��
T�Adj�H�әJ�25���?�����3f39=�=��wk��*�cO>) �AK��6
��-�RgƖmc�ee���xPj�i�ĲoK��ǊXFCS���%km�)� V�BW}�JmB�1 �	M����r�z����u��L�@l��}�n��]D0�{!S~�G��=j��R�pP����o�Y�x�b��0(��*�z�Og����(uJ4��Fzb�\����t�D��&a��Q0l�V�q�먴X����bL��q�����@�*P)q�~K+��ű�8����hu,�pρ�h�A�<�#��xZ-�a���?t�����)H��d/e#���������{Fd�x���<�����1�H� '���d@+�v�3S��^�~�US�T�Єo[G���A�����յ-���x�&�;���΍
\{S>��C��+���z,���Б2���c�Z]v�Ve��{jQ7)*M�3
�
.N2%��"�l7Y�[�̷�Zq��v�����~���y�Q���&u�����^Z�G�HZ�s}5�(�S�Iq�(�͍�����-?x��|��7Ǟ�j��+zh;( s��w��H��E�����V�?�!y��w�Bʚ�V����\a�c��@���eS�?|�}����29;��#�W��~���RY�Z�)?|�'r��%i���٭������m�A�=@1������R�V�A�� ���)��?��]����lD���}|鲬n�ǈ�펁f��>�&��d���#KEI�S��[��<=3k`��q�Ohf����/f��p꧛9?�+}��MF�?�S=?{�_����":D����e����=�x�\Tp�-����L�W\�[.i摝�チ��1���@]S��bM���%�G��Nm�/��g Y�%c�c�h��{x'}?�O ��ޒ�b��S*�G��ҋs��l�#!O�{9k;�eo8�(�)/����9v�Xf\Q�aZ̨�=p�Oa4,u���G��L��i3B4Ooٶ�e�ݙ/|��ЁU�g��'��p_~����%�����V-DrBiP��Ψz�A�
�ʉ��ͷ¡8T� 0����ن~/u ���L؈r߁jQzA;*�E��$�%����8�s#�C�_{�5u&E:A8V���c�$�*���(���&�p�}e�+8w6��xVG���*�9$�d���ސ��*�� ����b��l����w�T_�U?i���Z��TN\�/o-����?�������cy2���ML0��*</ bC�gT�JcE{֘�KL��ph)�&�����\�F�\`�E�o��dT�Dq^
���~��2 %@ڿ��rA^*c�z�%��m��/�,�������>$���UMLP]�x��,.�d�NSz�����܋���_���mߌ�!(
��w~�M���= ؝T�z�� 5��_�Z���)�3�i@�X�`��"]�
%6�CN� ��&������OZIP<|8�\B�%�;7��57�a�`�B�� D�u�DE�-mSQ�\��fc� d�������c�Au]:;��n����JC7����a�k�0l�u���������V�����Ѡ�sTf���n�PIH��5p@V�Å1�-h��V��jhKc�a�����+W�4E�F��F�B%ky�}�'��gݳj
藏�vB~�w�5V=[,Ɠ����}��q�&�x/)n`��G�p>᰼�uR�4H��_0H���^uDҤ�G?�P��ɩqr��y�~�I��s��[y���	΃O�e�{ĪQ�>*+�N��:���;�ƠM���k��SI�'��C��5Zps��n(��Ď:=����d��c�4��03/�����
Q� ��0��H|�pL��O�|rK�$���?R�wX�ϒ2(:��G�dDl�g|O�o�K�Ҽw�d�7u����#~.i��E�sѿ�9 b8�z�T'�X��hVyci�4�$t�jA�k�(o��Dy\�'+|����e�y���$t#��LؐYg!�����J����pq�W.]ޕ#��M��MWt0�RC���'�}���;����zĲ��)�2���72G�~�\�3�X
��q#�}k{�	3���&+�H�����L�3r TO�������:é1�2��U������)ߢ����߇�D�ē��<KJn�8t�H0���w���Q�m�yVY�Φ\g td��h/Wd}{G.^���f�ԍ�frC�$tU�>�L�7�2'::j�R��ܐ��$���n��s��AZj
Ձ['ԊЦ�ݨL�hR?-{5���!?~�]���~U�w�d{k]�9bŰ�1w��aV��<�^K�4i�q�����)���>4�b�
��-Uebf^�Q���nW�U�<�� �o����n��_�Z�2�V)szj��:��"f �q�%�������9pAq����%>��)�`�:h��-�;�U�k�55P�h�2%W�ݔ9���l�
��	T
C#�A	���9�T�P��F9K EӀ#�h�ixQ�0-���|<t���F/;��pP�Q�	2tT󮽝G�4�q��(l�S��թ�^b�=�F�z@�/�9�c9nP�2��ò^� .:�/�|Uķ
�4�J}����kC/���֙3qd�;6���}�ܚ	�峜O0|����(~��������k��0/�f���S�:N�������e�E��!�?T%=��"�){��z�Q�@��g�~J�V�I.�`��&*O
��@��#�yb�+�*˻�|/�X�1����{��ڔݺU�P>����Q��@��heD|�% �w�q��DqF�a�� ��Ĝ���"������wP�%�7d����2�fK#����	��g�p����0�<7�߾5�ɶ��>�p* ޗs��� x�kwy�p>9���:g4�W���L���	<^krk��k�<�j�����{�W~D�fG�t�R2��UV��MӍ�/
�0 d�^R�*[xy���f��wؤ�#��Ӡ�,�|u����iֆ��#�
��_2�M��Ir���h!X����%�1a� �#�'�0��k�`ۖ�BP*���~�!���7ΰ�K�} \��bu絟�n�����*����b�����7km����C�E������l�+Ʃ;�A���if��	�I"97
��
�x�� ,X�#�~zp��tWԷ��N��W���߾D ��]-J�Ǉ�'���ų�|���i���Vdcu��0{�?~\~��T����깙���	�C���o�戳�?t��k�7Aag=�_���*q��0IY��@����@h�L�\F�2CE�l��I[f&�H�ȓ���ՕM)#����C�Q��P&�K��`�fee]z+c`�<8��s.k>��c��7���2�#�еHIξ(���A��z���Җ3d��<D	���iP@�t�Y69���H��fCKU��Y[Y�'���p����$G��2�����ǕX�Rۭ��}���^�4�&�-	���a0�/�?�0l��<�'�,F���-C�qiR${߻������3�qN�"3���f�F�����޽��2K�"N�8a%�E�v��$��H�d�BHJCF�
$<)��M��ɴ�V�j�0�%��1�:/�V��ם��h�����+��33�,V��:�c�hH� �`��'��UBd[O��Ń��(�G�M݌�o�ҍ�.�7����R�Z:p�O������~���C�46/~�BPYfFl�ԁ��s�a�ZF��W[ݦͤ$8�$ր* ��sk�����l�t"�H����&�+�F���
�i^�ĥQ�Seud����J�~���xU��~)q��1־�2u2O��|$��P8SxY�9NX�
�������u��\  ���iJ;4�$�M:M����\�QP��b����n}]�'��H�?)+μ����%��h\9�,-gPN>��$ʯ���<�nP��"S�UMY8`�0��e�&�Y���JI��5���4b��0/im�A�����[wB�����*o���?Ca⨒�σ�_�O�l����O�Ft�7�wT���W��Զ�L�Nhp�H8:��7N��6o�V�l/\�y��b��{��n��ZܱUF�1؏��5~�sb��mG3�/n�?	k=��f�B�dPi7Ng�=d�@���r���z�~]�����PO��~�E�|vEm�H~��emi��a��ŭE��<�Z}=����^}S.�xRZ�e=_GzS":�<)M����,ц��z���vG��ZU M��~|T�sT���-g<F�`�lLdV�o����������D�u������.��?������>�C�<�N[>��3��y6���F	�I6��S��eA7��ڲ��o~�%�����ܹ��E�.����:*`����R!
5��$��e���w)�#�;�\�$O��9Y� p�0�il](�<�� ���q0'A(�8Z��a,#r/8}���T�m�q��AG��ǍT�g��0�\�,�)S�~�Z�T�O.��|8�q\�7�yn8��ڡ���8�9+E�pc=r�*�y>��8��vf�ˍ��a�'%4��x�|�_�qoБ�G�j��t.��{In� 8��N�z$�2&ò�s̙�fq��ȁ%߹w[�ܿg��Ч�T�DH娔a`���B�sb:D@`�Y�_$<|�`/B`���Fִ��o��!De��������o�HT��)f���ϩn~�q=�8p �{-�2�(eex`(�u�v�$�qx}��-�����y>p�Y�7g���e*�5Z�+�(>D��F>�����rf8�g>���ͳ�;C�1H�؛�TH!U%TYuS"1�'P��>HE ��%ځ�q�W�I��(<2�#�?��ZNu�٪������R3�p.U<�o*??�B���g�FZy����TXnU��4;��	��$4AE����VQ�Nt5��x:��:w��c�����t���@䧓]X��&ӌA�F�`gq��fW�.e���{anh� �՚dsK:�pl�HS�y�s���F,�}����oߗ��=�77��}r�R����<�����O?EgH��;������2u��V�q���n\�Q��ǒ�Ԑ��?�[I�1�8 �z�EYo��Q)�_1�FҲ��}l�=��S�H� �� jL)\ѩ���zm9�U]W/���֞�xO.�Y��f&���xp.�DPO#��-گ�6��y��4����`O������wi�����F$����F�tj0u�2^>8 +�	^��c1EI�����P�M��:i�D��`"�E�:A��t@z��;\��Q�oU�0��6L܈j�q\
%5��*~�C^�BE�Gr�(����)'��߇;>޸k�j��3�(�6>3K�SV�`�aXО��
����d�g-��B��Ǭ�k��)GM~�ړ�騀\��.Ķ6ܗ3���"��xL�B�H=�1��	�iM�05�����C��� ..��'FƗ�W�'#�VT�D�I����HB���:�h�?������p��ڃ)���3�0�C�'���2����"�H�! �k�!��d������,�p���%�i(7��J�&����.��p�Y��'��Z��������o��8�P%�� 6q�4�H}R�Ӹ&\�r>�*�)���~��$��}���熷"�3�C��ʻc�4i)�4�3����y�������t"��Ç�r�{(�=�/���?׈�:���܏Ɠ �gj�$)KE:�'��Ն(.E�$�lR�M����M"��-��,��qH�93H.
�I�r�j�W_}�=�z��;" �c�S�ᥗ�Np�z�倘8	�g��'�[0�:�ct�F�P]?@�6n�琈��a� �HLLé��Tv�(�Y[2�8O3
�P�0 %�� R����>wR\賀�����a�U�5ה��5i-m���!����	w��:MV�\\_�1CSP8/'�#V�w�8�NoC��\�3�R�`�	�����|b?!)��ixNS�-��T���9*�>�2��`-.�$b��P;�ܐ	LHL&6��$�R��y���W��ټ���^3�'��.�}�	A��C'��d
h[�N������K���a��
&��A�<�Z��!=b�+��\�0
ʎ��?��M�0.�������@3�1%�hB��hO`�9A��Ĝ#h8��|:T
�3l W�*�
=���E���L�'I�<^��N2�$�"6+ITyC;F,�*�}d��?��y
�<ꦄz�X����q�S��NX�~��6�E����������:-��DRK�I�)��u��'v{o����k�;<ܥ��S	G-�^��FmL'�48!�G�N �(b�5~�~��)D���]���h<������Y�EՏF�*���ylX1�Z�U�3z��e¨i���H�~�]�������L� ���8F����z��re��Fĉ��2uqK�֌9���L��H8��SG��VQ��ۺ�J��1{d��L@�vЍ\��q|��p.0'p`Ф3Ѡi�a�I�
)��Uϳ�'՚)�r�2��1Aa�����R,�@���k�i��t��Ǵ-������A
/p�|\ �G�JϡՁs}|��϶�I��?�C����u���,�پ{�x�05I���׃cU�Ϲ���F0�A� 	 ����U�"/�v{�Q�}��ڐ�5���(3]5
s��/F�C[��k���&Q���ž��Zg��`)���;:&G�>��"4�,,�~W�lɑ:@�!�*��N�sHy��QvJ;�2v�p�hၯ���9[7&I�!�����<%ɶ�=�E9�I�䃷.G��5�[��Q_��<����X����C9N�`��i{Oע�G=uP�/?)n|F�fO&I�&ʜA&G��ĶK��="}&5y| ���1�s4bH�`&Y<����[��f��	%�%V�ee뙳�����D�z���׾"�ϭ�ރ�t��:.[�r��������-���|K^{�MYYZ�����Յ�c>��;�VU�8i���ƌ���I�s#� �gX�!�I�։�Ҡ-7O�Nhk4	QuN]�8�d�(����,G�㈕�y3�i-�sZ��&����"��
��"��:M�S�::=
��:`�{�	�*�(��6�:k�a�G�C��`��O�w��Q�V����!�:a���;*3F�����~�TO��쟔 x�H��Yc�S��G�d���5Q<!�(N[�{���$������[wn��D�._�B�KQ>=�7�L��l}�k�k�II�<�"9T��Qe6�Սe��O�_?�(�vi���:�N�8Dl8QG&�t��M�fp<j�^�f�M��@����.��P>ϲV:�)��,@�qY�&1KJ����ҒfP�hj�(�A?��0����	�:�Wk�,O�U��QQr��a�C8�ؗV{L��ѓ|�@,Z� ����7,��ۜ��ȅ�m��Qŵ�P�h�Yo�� y�Q�L�7��T~n�I��A$ :��SJ��$�jLz@Wh/ĺ>G��B�$n��/�=w�;,>`�:����M9��E�?���81��c�C�3�yY9�t�6;	B����ϭ�<I	�Hi��D�8OI�G���cOƵ&1�|�]��v�URH��lW��)SX�@1M�L(�h�a�h"�m�3�DD��0㪁�[o�%W/]�F���2�u�S4��T�Nʔ��������4�ߍp���Qw,�j��3R@PE��s���ugFf"�F\�_,2���Á�X$���\3�Jk��\}:����n�a�w0=��{������	��LN��h�g����Y�]8/�g/K��e�����3y����D�ѡ�U��g�"���"�	��B�yA/�M�N�9W��_��V@�h�1R=El"K�rk e��k�"˿�Q����p�Z���w���g���������SO�CT�s�/Wn<)�V�,��X��� .��/s��1��]�m���
���u�b�:!�Q����)��#�+���B���"��"��F(��C��J�@�	��Kكb�Egf:6u떛V��j*3��������c�g:����4w�6:b�����mNRn3V,}>��*����\D����w�%rR����+����N�@��Q���?#�:�2���z��r�=��w?x!������?RhQ��;I�arg��	��w�}y�W��7�+�+� ;c<_z��|��ߦ�	N+80��0
ʲR��4L+jt���+��)S<�����o���{�C���Y*���(!k��2�qqbl�Qy��PL����"h!���D�����g	�������ĕ����3T��\�ȝ�y~�,��q.<-*���˙��Vq�����Q�XK'9 ^S_�E�V��
�!�e��WT9d�ذD�k�kJ'��&�nn�`��CD�68�1��^�A��"z'<<ъ�uh��B���}`^�HN�Ȱn��Q�mX�����s����<{�v��
��3������_�W�-S�b)�8�ħ��+2;�eb}e�1����Gm
.V�E�83d;����I�Dj3S�I8��Q��#�.7A8T�d>���Y5�s���'�g%l��>
��������b�((а�Y*���I�T��!G��C!�X�Ԗ:9ݍKr�9�^�Ý{���8��D��<ay?��R��Vo\��s�d��5i-��(W�G�~�#Vq��c��Zf$%JU�ִ�%��������qT��H�f�u�XT�|d剶��*N�hY��`�
�D���W_[�����SOF�x�I�h����{p�Y��nu��h1��(�3]���������ݐ�A2UNka�U�?�Ԅ�+I�yM���i��bʱGU�gJ\G=K�Pi2������51 ��:�䜕6�����i�)���V.��Ă�M*�ϡt�U�����
�(]���D���2���@Yk��Qi0��w�ܸ{�o	$c�W���~��F�RT��LJ(�CloF}�(�\���}t�{��FD�B`��=V����,�L���QGd�L��0p��)����	�O~�9�.��ַdi�G�:*�����zӈ��o%�g7��]��y(�^�I4NRKF�B}8_��OO�0Ft�8G����+���P
�blMӲܜ`kX��mR���b��6���!1����1��J_�U�ߏ���!eکQ�]��dsaQ���7�.�������c2��<	���YB��sg|���r��ç�w�������y,�����.��t�[t��Q�-��m�L)�kYʎ���Ȭ4*�����C"~���}�>_��n��y� ��Du?$� (�糈�?�<Z]����tH�g͖!'�?���`p [F���enݬ�"*	ɨ"euXҪ��*���@xG �h2�5�=|����O�c�I��|KQ턒�Ԑb(̂L
N,=FԪ�Ϳj�fN����&A��9�f������R���eJ���Uj��{���t{��Y���\����p�Td�<a��u�g�i0ߑL��d��.�"awz�v�,���퉓�����4���d޺$h�`x�~|L�sTrZ���󔇲�L��(�a��=�,�BW�"T�D!wQ�F�X��W_{Sn<���7��ӟ�\6w���kl�a�ڀg0)��}8��z�Ӭ2rDw�h�4�ER�%2w��?�X����'���(ƌj��d�E���H�%��a���6@R@����N-��@��X��B�2/��ȕ}����I]��p��Vz�$|b� �mn}D #uz2$5�de4�
�^���BHf��y_'�����u�"��U��?����F��0��:"ue-F�88��%Y\^2����޻f�TI����^P�6���Ҳ����f�Zh�esut|$-5P@>������������Xd����m�!�y0r�P�Zm��ޔ���oB��餑�Bޖ��i�h��q�D�|�S*�aƇ�(���?Bs��L&U���(8^D�J�3h�p�*���n�\���/��dZio���}�YZۈK>���:����ȟ��׊�����4hXyg!��8�<8L����S�Y��2��E������r^ʟ��+��C��dsڷ 	�7�5��!��U�a�H���	_W/NB��:?�֒��G�<B���������_J@�c��#�LQ�Fx�N �bM-����ܑ$O�(;�Z�M��<�@p�:D�g���B��y���n��ꊴ5 9h�qt� �T����26��k�$�ɰh�G��Rsz�qqBr�Ec`QHq�׉D���2zށwYL����M�5�D��#�F����:贗eq�#gB��s�B�9�� �����Q�8�/�;�6��a���YKh�Ĵf��8I�^��O=���o��#��P�,�v�?#��*s�Ib��#q���F
�`8B@؆�B��ko�#_���ew'���������`��G�Hӟ����o2�A��I_����*"��U��U	mGqY�-F,EHeE�X��I`Vދ�!W@Ȱpfpa��Ό{+��9pw'�L� �Bo�ߛ�&9>��sqՕ
���.���n�� �fC���z�#-UAF�ī.���T���vC���S�J�CfS^��BR{���ؿ�O2�Y`BJ����#�(����d���.�y؃��������sCQTzꞒ`0���]�214T�P�#
c��~6�Fr��-������-W�^��gγe:K��gON�y�]�Y�����;�ģ�6o��z$��1*v`$���i q�?��eѰ�^�J���br��;�T�U<`�:M�K�����wRA�q��x1��:��/G�\�+O�%�ڝ+!"'
YF�y�; .�����除m�Zdo���r��&��;M+)�r�z��������)k;
B�� ��V]Oe~q�"D�q?�#����qj]�4K����r��l޻/�Q�6nI�9�zp��i����#��rB'���H�p�8�1��i�`����W�Q����I���g�,�uy���h͊��ܔ����q.�����ɑ�4��#�"^��:��?Ӆ/y4EQ9�|Ӡ`m�|8�̞u��Rs
��jv�h��Xn߿'��o�rr�&r��v7p���LI��|3`7*;�U��>Y�$l?�)����'�T�(갂X�lY`��L�_�m��|;&,q�@K�2(�m/�F�1�t��V��F7�%�G��Bn�ҙdw�ڌ)T �)1˞tf���N⣏�|r�iQL&�x5h@����Y���q͔3&����i�C<8�01�ҐW�|O��B"����9� ��hr2�0� �C=�I��0R��GH�2�X�M�>S6E�'���_���Ȋ���S�x&�P�bg#%Y��(7<=!�Ȧe� �`�y�����RiHq ���Κ�5�Q�F� �Y�43^��Ku��Y:w ������d�7B� ����}6&���'9��Br-�d��mȚ�T��\Zh&�#2cH�N��<�owp�X��ѐ���	���^����+��i�&o��˿	�Fii��N��/PUet���o\VG�:�U&v�
B{Л�[����tخ_���X�ݸH� �"BI R<�Uu���v�tF�.�N�u��$ڞ@"3�l@����W��p2��	f�"���f*'��+��H.���E�@4M$)K���I���C�bj�sf���1�*�<�U�KM�F^Ε���4�J�8�S���~�:pIw6=L=�F�}j�\�t���2\p�`�A��z�{����V��3�I�lTk7/�3W���|��#�0�>.��}8�kk�����K��z��+�����é���`GQ)dÌvq��(lF��q��y�MC9V�ׂ&I��8��f�qZ�7�(�e�0�ߝ妔HA!3�~�ɭ������ː���,���I[�X����ζ�������_��q�F�HB��1�'}�vY�b��f��ֲ!���y�(��l�F�,6�d��ZE��X�i��#ˁGPL-���C�G��w�ꬤ�~�3�Ee)Z2,H{a����c�����F��$��F�Ƌ��3�Ÿ��,�X��s;���)ԠO7�#$�)�m㾏�g�az(���4W#9%Ŭ��l�4$8!%W#���j{�Ly�Y�!1�p�������=�ڑ�����,/~<���<�/�	�d�Z�?0£F�`���>5A�bKE%�lܶ���ΦE̼�9�QEd�]�>�=	;B7�J����{�7��M#1�v�?1h�eD�cuDX�܈�U�
D���
*�d���Q����4X�[�א�*2�ã�����-�,ȿ���1�I
�,2:>F�Ltd]��#�T�2�<�:�ü�Y�	���sGu��"7���\�!1a{vFI:^we����-��0?�L�&̧�1+�����5[�C�Y��Nh1V ��cD$�0g0&���P_���$���ѡ����tr�)��F����z\��{ƪs�!
�X탵XD&�>�C�G�U��ro�$a��#�e�C|lM���>y����O.:É������:Nd���~䓚�[�28�V	f
�-��npw�D%��A:������۴�eT:gY�v��fA�/��xW.|c�z���~C������ɟ�����Q��4��%D�Q���$T6	�L����
��N_��T��w� �;��4S�����T�Ϋ�����;��a��}�����JT�ᾟ������K_�"9��;���yC'm8*��9w��~�qp,Y�q����~`�y���RB~��;u�,̭9+��O}<�)h��%��_�J�6t6�����/�Ē�w�~��*.��&`��㝼��y�v�M#ih< ���#K#��B	}=WPz��yh��B{b\8�}�,.�&އ�pCj���R�����+����E��(�;����"�#�����Y��k�ҢړH>?�^ 		Ǭ��e�(+h�[�pbǴq�����O����6��U���2�-�	�b,"14s��G�tO���Mr�v�K�lq��
��p�W�(t�!��<;H_�%�߂��wx��8�z`��e�'��j�92؀���9�p�AԱ��u������1
7�J�Xz��!�|f��[n���`T	�(�)�8{�&?����4"Q��#�X����UFop���ٜ�>�� P��j���K��&������rS�9$mB^D�ݳ܄��a����$��~�@ѐ0g�m���Iw�WB�xJ��{�-��{�8����:j�G�~��<���L+�CU=N��D�K�}S�� 6	1��H>"��F*!�n$��������.^�&�5����&}�xP������N��r�t����OIrDy��K�v��h�u�E���,- 
6�J������rf�'+�=���{a���ꊥuot�~����⹳��>'O~�Ӝ��߿�6o���������m5��)�L[�F�Qe�9_QE������k�M��ˌ���1yR��#����I�n�P�L<п��/�9�������L�J��$����gF�&Є��_'^����׫Dc��A��n���xNj:q_l"��M&��>��(�|��1��̳�[��[�nN�l[p��=y�wx�������pf������'�K����O}_=:���Y�e�=�_�m@�� ��կ�@{�]Z�����F��Qb�)B1sIo���@[&��D �O��v����u��t`��w,�Z$�7��4�-��88�%#U��b�� �[�1�?ݞ�ޤ@UN}��E�v- �O��La�&ƻJ,x�g@=v�����*��(��|��g";.�FM*�T�ۨH��z6M�6�pW�\���62��f�؂A}- ��tG��;*�f�A%�P�c���5���U C塚��r�c���B�m����Ӈ��F��%d`0��� �	@	��4B��89ȭ��xI����t�-p���v��7����^�7��F�����ia�*���̧�F~������z����Q�&�v����p<F��a���c��/�}�,w���L�ܾ)��<�Ob���Ů�Ji��:a��FEB#;,���8ABGV6���3g�F�޼���:��ulN�k�$��sGK\~���G�k�p^�lC[[ݠу(�9��d��;IR�3c�����#)�v�~��n��~�a}�p�|
G��&���p*�%��݁�q��k�8��0�*�
	��ah�{	��.�52�;�r���l'�}2��Ȃ1��8 X/qP�<�H�ЗfC�����\���u*�n޺e�!��5���Ԫ�����O]���o[e��Ձ�1�'���b􃃉cδB��m�u�Agc���NIR�wX˹Gq���f��z����ݑ�;1��Nf�a(I�tΊ����L*@*eZ�1O�ʥc�ζz���t�X���H=��G��c�,TO��NL˂����9.�U��ؚ��u�ϙ��d���u��G�.|,���|q�C��S1`r��}��36�(��>�G�Dm��Vdpz,Mu��?�GG���3t�<Ѐ���5����b�D�vkE�S2Zԛʳ٦�>�>V���f ǏC`�J�Q��{v���zq[Q<2>��UO�M�z���^��{_/�3��f�*Ĝi����K#d��qv`[C�#�����?WW�I����m�c�{�����i8ĺ��=�u@UI�Z���$fs���̋(8�5KL,��*m�2%
�FXc�I�	��`m�� j�a �2al�NC�
�'�	�RL���*����L8��VN��,�B/�l�؄NRs�ω��yUϸ"�T85�F�1QV������C�Ŀ�� �v��7Zr؟����Z�;Ǆ��*�a��5<�����￨1��70'L���b8��T��'��Dv6w�P���������i.�A"R=U���ugd�C�E�?������D
����)�%H NB+�<��<ڤ2j��_�vک�������Rr��3:>���������`�Ɉ�Xį��������w����}�,���瞓W_{���4��3�yG,]�Ј�~�4g�G�E�$W��\���}������bΙp���Qup͊����>�0NJ�`y�.5Yj,1�5BGO�����3��'e�s^��Ȍ)[u�5�W1��,
P8����Q����r�Q�ƙ?�a���bs�&�EEp������&��Il��U�)$G���Ɗ�s�/sO�����jw�t���?9<$�"�ݝ-�;mV>����8Cy�����ӧP��߷�&���B�9?ӊ����D�?Ƒ�4�$�+�h��i�zT*Q�Ga
��u�iDa��EM��׸�Ӳ4�=����St-1����5�����;t�	�B�y�k�sX
�4���ӂ�x^\����k����hӼL�䁉JR�a�+�P��6�p�9�N��BE�k�TD�l�9.��ʼ,�?��y�xQ��6�V��_ދJ|�G��e�ʊ�
(�{�y�[r����~�V}�S�b���S+����$�!n{]"6"��C��Il��Í��iE+�e�J��;>��#:@|��%]�	�e��A��>H����}��c4�]�"<,��M:3�A� ������1P	2NM�.7fc��DuC���x����F��c=x#=��egT��Ћ��Q�D'����u2�Od�?�I'����,��\�G<Tq��Q�B���:2}vI�Bd���pp*��O��h��C���ɐek�dA	6џ5�TDl���@��p��ם��!�B#*��nT���J�`ԫӵ-ܧ:8m|���������|�/˓O\�k��k4ؐ��>��3���˫����'?}Y~����� �;�s:5���3�K���4OrtZ	˾��5��Y~��,���ZX��@q� ����񌑇�.#)fġ$�n�J�jQ�r��:W�~>�p��{��,��)��4��'�Crr�pOQ�v��ۙ����E���g�^��F�1=	��cýZ��\�\Y��_�a�I�-{�8����vV>��S�j[�]45�[�(�duN�BY-��l Gs�z8X��1.���d�i���U~���������{a���4-�������h>O��S:�sF���YD�鄪��ha̤"iZ�]�b�!h_�A���Ԁ��"]'����{@^N�SF�%�[[w�{���b�;kq힣�e�>���2oQ(-�#V6I-e��+ �9n��m������w���k�jǆ(ƭ�Թ�)���QN~$�n8�������[a�*��;���d�Ҵ�m�P��_�:qoz�&7�ˤ&"�z�vp�烢"�).G:��*�?HwW�蜬�=ǽ�f)���.���[�	s��e�@(�_�`��𣺧�C1�'�sP�p��m�z`�%�g�[��>����c �N��&�b�f@&��_�>dhj{zx�T�ѐ�,�k�Y�����H���ak��!�[���O�]�lؚ��Ŵ���V
=㢞|��#��E�m7��x�����?&I�l��D�Np6����FC���C^�"h-��MH�,k2�E\<�m��P�l�Sp:B*&�5�'���tA��X��C哝�}�p�Cv41)�Ӂt��%� �z�8����h�d]���� �38<P�-B�a�h�������:�%��}�y�����_yANN����dmuI�ѩ�.ˍkW$}��XcE*q^�º{;a�B�����P�8�;���X3#�ف��W������
 ���2��U�y��C��:!/	��;���3L��$�)SD��9�?��"14�Τ�J�48&�m�q�b�5J�m�ib�0����p�*�[��i)�x�,�ĭ�mD̈�	�keuCΞ�$gϞ��9M�wo�{�ߖ8Zp�aLp��P�Ӳ.�xN8�8��:�E�̩�w�-�<��Z�h���Rt|~5爖l��3GF`ƹ���g����F�N�GR�>D���k�VJ�޹��>������{���@�(�k�E-�ܧ2
�r�����k�r�%��~���#�U
�D7�#��	�b���w��hWzܬO �c�gK��������~��pPp��N���"7eWC�;��Q�WH�T���:J�?�^^6���d2�4���a��X��/���d�6��G�95(�8�U�EE�j���o 2@Ϳ�L�П9{�h�h�YʇI��:���ݨi\�B�K�`'�8����P]R.Ediҏ�0���ġ8�NuR��=Q�͡�]�{^*Qy�2 C���g��z�,-霭�r�v�u��0d�||�P�#9��)��0�݅&�z:R����f�ѫ�؝~Ѥ׮O�QY�,L�\:?i���ڒ㣑��i.�d0���V� *��dćM�|}�R��@ 0�#s`�: `+Ce4fI��T���[!n�i�d�Ѝ�|`+H���K��d����|m�O��5d�P�qߺKb��[���̯іb�R&i��,���|��z>L�}bz�z��5R=�c��CkYJ[_&��r�ܒ>K�Odw����w���u��7U�_��*� ����%�ޗoh�@�h`��Q�$l��갽�q�7��v���mx�:///�3�<#�>��ܼy�<�)-6Vp�ʍ�QeZ\u�E��.���zT^ߌ~���;�%�.��p�/#>!`�0 0c��0�,���9��6Sd�<	�s���^>'/2������ٹ�4�]�9#d
��}.!R6����9���1À<|�%����{A��h�ds\�n���{� f
�0��82����8%���1QD�#�fk�����DdaC{���NE@�����jm��s9��QY4�K��E��e���DN�ˬ��|o�l��Lm�����+�P��ô���|�)�� �njy8�!U�@.9�>���vx>���	Ε#|�Ly��)?��y��6����PmH��jP�'��t6�P@�YIX�ޅs�Y؅;�r?�E�h�~���B2���c\��0D�v�3�G}�,�όC��̻u>��AG�Y��068d�����9ρ��灷������_ѵ�*�C����7=ʚm�����8�ì(�Y1&� N�K������j}J{��]����Ď��)� ��G��j��q:[�ؾȩ��"7p �H遼��FZgX��z����&q̴�+�색�� �h|*�� Z	Ni�
Е��Z*����G�ǿ>1Ge��̯߸����'tP�L�V�ey�lF;�w�g#5� ��L�bOՐ��iA�}Sm'��-�k6M<���d��hj���\���]
@��)p/�"��]������#���l�Ut}���t�|���
�|���0h�!����|,��#����|L���i�\�X���`r�t��I_s��#gϬʅ���@e˯���|�3�����;ܒ��5���TS#ʖ��d��A/�8$xv,Fb���(�G.\<'����L���/����C�y�@^x����u��C��?��;.���j����T�_���z���}�z�3g�I�C����g�O�w��]����+���"�����Z^�ݭLĻ�2�f�k`g��������5��e��)5b} ‖Kga1�Z3�8�!�+�4��K����g�ݺ�s�Է �3��t����;r�D'ԡx����}*�r�$4nl��}O��H.�����S�F�y����i����k��Ed��:�{3;���F��)Qs��ב=G=��G��r�~���%R���W��L��s��TL���VxI������GƬ�³��N@XP���V__�F=$�gw��v�s`�NK�H=�ɿ�T���xT!Ou�r��ѽY!�Ȫ��r�
�5K�y��Ǉ��㿏�M��v¿ٻ�Zʉ�ƦA+�*�5ܽ� ^�Al���� ]A�Ip��D$��o�'��ps[F���Q�5j(�������k��ǡpQQ��2x�Jch4��.�8K�p	z}�X��[:�}�a�����G�x���B�˔{y����ޓ�VO�l��{"��ѧ(��-^ckMU_-��!%�ިͤg/��>Xٔd������
�R;�3�����xc���u:zl�=�9bIq�Z���i�'��Wo�c�㐄G+�f'�Ɛ�AWF�ly���;��!z�h���X����H?�(�bY_Y�C��Q�dz[��q/`Y��!R#���`3Byi˼Ep
&Gt�D�u6�/L�Ȟ��iPXYr����=�y��AM%�x-:�brѱ��r��D�8�t�tne�RTU�M��L�61/���h��_����������5��{ߠ�ƽ{����?�PV�Q7��g^�®ztc@%�UGL�U@�g��K�̦�l{l~N�'��*+k+���$O=�$��_��<��S���^�D���K���A��^�R�Î�du���6�R�������ف`=���A�fy:>Z��d��������]��}�sT��T̆:)kz��E7���0�j M���.u�Q�������e�QA�h�F�u8��V �=��I��©�Q�fL��9���K�CF�'��\�RU�ؚ���AS",q���������J|=�$}<f�B�R��A�0�,p� 7 c��I����MQ��"���P�{.����F���!�G��[˅8j��︣b�]��Q�%U\X��pf��#+�xcp�pp�C���&wp�E�e��:���ޢ�*�T�U'��A@�K�uv���k��;�Ϳ�>dx��TK�(��V��PO!2��(qD'Oz�$�L�E��A�?�a}��'e��{[�e��#��q-��Z�=�-xg�0˸Z����A�U 0��H-/1$U�ldiEY�  �#u4�,v��k�8��v�)[O��࡞�}V�`�G�g��.�qW�<)m�W�d���{7n�IdB�������α::- �	��"���T���ܚ%��?����'%�DӃb:�6��yvmU�X#���	E���!�Ɨ�W(V�����'C�t�K��մ�-V׌�
��H�d�Z��"ш*}��>�I�i���.�φ�'�����0�ۦ���9������<.P~<"O�]���9�aBI6UO�>0ؘ@x�
�u�́p���*9F��bS��=m�uXF��G��i� JU��,.�r��F0D�(G)2x<�����;�Hی,ro���a���P26$�PTǌ}�I�ՕS˯���ݢ����y'�y4�uPܐ̓���#Q�|tt�g  (RE���ӂ�Ƭ��b�c8��z�c�Q��	|�^.U��T���lnP� i��t���<��0xG���i�,'�G�e��R����p�FbQ�޸�q���|�����wx��ф�#y'�Ѕ;c�,�|���h_��"�H��NCX�Z��(Ҽ_�7h����K��?':�R�������l��:�u'���î(�eؔE����Q5�F� B{Yn��U�E����>��Q�4�=�&���Pܝ�!�P�<�4r��)��4�0�^�T�tc��\��⍀���s.#��i�U�Zwv�wT�?�F�>��}8��|�؏"4��^@|�54A[Z,Y(�@�,X��s4x�����D>	��^±�}0_]�FFx��g�˱��k>-��'���~�n�ӊ/���D�x�	+V�1�k��� �$�q�bܠ��4a��P}��m�p���A����0�#S?��)&2*9C/M��|0�QhlP~f�^j`��}��Ԅ��"'������ȥ�w,{[��}�=9޾�g���}���瞖k׮ȭ;���;rs�n�աh���+r��S�i.e�S���>K�H�lǐzg,�@2<O������9ƀ m���Qi��O�a;��8��D�����eX��H`xV��Xv�M��Q8d�4J��a<�H�C$�W@jK�:;���F�X@�m4�A^_r8,M}���ړ��-IԺ�T$����Ή�nX��&������M���#�-�R��fʞ=);Vj$�Ad]4�M�Fr���s�h���{��h����F�CY�.���!��!q���&�Gc��a3"��A
��<.̃(јݦ�Tz�&Y� ��L-��#R:&�oD��N�l,��'e��1FH���5��	�d,-�Δ!�2�q#ب����J�/0��̬�؜ :�b������E`���Ҋ)��F8^�()�M4<�����X$_��j�����BIj&��#
c:2؜�K�ѹ�m��g�렷�$G����3 �)��k�j����ߑ�>x���
��NdKt���	�����	�K@�(�<��v��+��Cu�A���`��k�&"T|��A�xw�P��4"?Q�-
}� 1�`: X�.E8t�9Y� B��/�ЭJSC����S���� -E� Zn��i��=r���;�S"|S���u��/��S�)�y9�?��D�6�v� 
~�*^�]���%����yJäb:���؞χ��y0��σ�TmCX���@Ɓ���=�/�%�%��������Ǯ��S����n˚�Qcc2
��U���>T1zU���Dc�u:ݞ�}G���C�sGCM�9.	��1�?�S��0�5,�Bʩ*K�:a���:�t�>:���3uSwx����Y���-��{7? �������	��v�߇֔����Q ó0!.�ϩ�O�m�N"V��8"�4e� ����H���[1�y&��m8P@)��hK�ZHJ�ǀʘ�����FW1�E�Ӂ�lj�������I"Q!L���8�]���o���H'��IU�z+�]�(�z���-.Gr����M��O^���$��ʙ�O���s2���>�_l�X�<Z����ň�:�Ŕ���qnJ��x��(Y�epT|f�puq1;7�%��A� YVB�*�ђ�n�Nˈ��F�V��S�|XWJ�g�d�JG�V��c}�)�X���Ҡc�1kː�4���� NGĮ�!�#K��CrGn&�!d!b�-RO�=���D*���Q8�0�����&Zq�id֖/�w�lm���Sש�	b��˗demU�ܻ+�zx�b]N��b'NMТ�	��:<�i����43���#x�Jǡή�U7�.	�ʴY �����g��zz̟a����k+8.Q0�P�8�غSpM�P,59��{~nG��[�Q��t*��-�nD���p���6����?ъcK��g�����=�i4�j�IF���[zkp
���/_�+ׯ�����lnn���6}]3���vw�����rT��?�0!R�X_�kK�p���p����?x����������~��?R{��.�%����riuE��P�)q�Cg�eb�[���S�#�f�0Ķ~,�F�A�E@��ta?`�`|�p=I�8��!�z�}��	_ �wߑ����{ ��xk��O�F�%w*��3GDb+Cwg���|kH�eZ���I�����*5�v�T�-p��و� eHa�bB�d;���@���c�Ux� ��g;>ܗw�~Ov6���W��y_�,�kՃ�p�3�( ��t���� ���yE�G#�u>ۣ�U�dk
��߿/������>�3���+��S;5�������2�Vi�оFF�f�b(�F�I°��8�`��=�3��lF�z�4J8U劀㞆3%�f�	{<��o0�d2�;эJ�{-�E=7��Ç[�w���{K�;��Nd�	U܉�]_a��=q]�=�-�w?��/�W��Yy��we�e�)w�}C�w�����eM��%��E�3������:G �*��3�*�h����:*E�Q���'�p=���B���{Z�ɉT��m�я�z O��+#��J�Ĝ��8i���O'����V�Yd��&N�c��P.�>"�)���$�!o���POݰ45�Rh,���8���r̆}I�ʬN�D�l����
�R�2mK�����]h�ʦ�m˭nRh��`�T���챡Z�"�����w�B0nx�����΋�ݩ$���C��?r�F0俋Z�ؚ���Ծ_'��r�Ȍ�$J��c�nV�֯y��\Wu��yF�qe��|xTKuD��YH��!jQo0^0�X�W%��f������ybe�ʪi��;5	
�E����şB�!]A��h c_�H~5� F}Y�=����>?�W���Yo����MM��`�p�ǳ�g���-:�7o�$Oc����S�&�99s��HS��F�'�o�5VP�;��GwN|��Q	���_�,��<݃�#"G7_K�K¶;�����m)���(c/�y,�1bF��)��~�󸹹mU�p��fHET�`�"8B$�a�8��������ri�.�=�ڦe�q&9N�S���4��>�ҍ(�L��[���$��6�OC�������{��;�����z����rR�����W��	�6)�{C3�]L����*=/9�-'��7��R�7x���)��<@�1wX/���s���ް�\e���q)���̝����e���_
6�m�!q�  ��u�`-R�(.L}٥ȑkv�`���u�(��Qa�g��B��-�\��E�HC�]Y�]y����`�N�PV6e�y��<��3��ӟ���5:D�����k�~fCVV���`���kwe[hT�fI[Zk�q����B�CL���'�_�K�Df��������iq�����^�(��[��!�c��U���Hbvj��36<��ŋ�*�����epz(����; ����X�H#k�K��6zm�[:�,�=ψ���a��n�װ&�q	/��Rsj�>,�$��y1�ԕm�[��{����Ң�x�H��ŋ�%��v��9�u���G?��|��+���fy��H3�=�� w`��f�]�]#�e�pL2;!�\"���r�:���I�����,�J��i��Cb�a�w�d������<�`Q�BB�<|?�	w9t����ipL$<�WDQE��5��M�xͅ���1��'4�pT�W��gq�2��l�?���L�FhcK���F'k4������2�Xb�4��H^[Z�t*����n�Z�<U�rޭ�Ǿ����Q��e����H;Iy�q��t<��*��2
��GT*�l<�C���׼����
���l�H+��~�}� � �!Cj�o�G}�B�Y�%�V��[#!�/��I�0��Uh�(��/���wn$�r̈́����lŌ���̣�QN�<��ш�9���"�IK�E�c����S7RH#�L��>�78*�Z�)��� ��Bs����qU}�������ߏ���ǤnJ���k{���t�yf��Va��Z�1;G���������Ua*�5���I9^䦕�o�`�;y:�N�k�$X
}�"�z��>�ӑI�?xe���,y@���jS��{-9�ے���!��w5���

����/��_��\� ���o�u}9��x�*�[0�K�/��K���]Y�`l����֖�Jޓ��YI�=A��#T�f����Мo�ϸ�A,��-��E�9��H�h=4J�8OB�D�6�3�-ׇ�b��B�"K�M��t���}�_����-c=���n,F�m�p����.��^���3�C�J��{�Ӻ�[bS,M쐏M�� Zd�d�.��[DI՗��f��m"��j߫+��^�z>	���z�(��A�K�G$���FC�����`kO�V7dqyI�V�������^L
�`�y;1#��~7;��U��3��I'�|�R�ud�ŋo8�\��=sa�y���;��{�g}�<���u�M���0pb��i����31�V��,:�\��Oh�gZj�{����� ����s�
t�x �$ !\Ѝ?m���.��`(���I�����US���9�|,t�O�{�����)B�f6뇂(��{���P՜�?78�az����AgS3�K	�㮝jw⬧,q/.(�����z��;;���}��c�J�OG$6�M@��aO�fx:�9��NU�\�=f���<|U�٪�}�d\	�Q���a[wP�um��b���ًÁ�/u.I#�K^��a�b*���[f��Y�2���t�eI���{�5�aW���*�@CŌ<;�*�q����1��;)�6�K諱pd���Y�� =�|�} �&g��-R��Dl�Z��ۗ��HMy��Z�������Z@���)(c����Y��g�CM�>u�=D�"0�a������ͅ��;MYꤲy�%�[�I3Y;�,�V��xo�
��/��z8�w�?��L���'�qv��~��H��p����ߡ:H��~ ����M9{iQ��NM�9v�MKYeW9��\� 屳n?���9*-�D�D�ż�Qs�%���@l�����X�I��$!B�<���|��[��}_gW ���oi������|����ݼ)g�^�s�˥kOI��Lh=%Jke��� ��*�`��š��bc�7peR�X`�ِ��2�w�]�"7#�D��7P8 �G��t"��;���]���ܽO��yh=�ޗ�s�%jvHC.A=_k]m��h'�5�
Pz��������ۖW�>�^sN�L>F)�)=��kRy2)����5�X?�~��2�y�0�X3/�A܋_jFx2�|�N�l��h�B3"���g�����X��k׮ɕ+Wԙ\����˖:3���ț��Fdm�\�D��h�^H�i �<�K/�$�ԩm����M�9&)�$n�L��1CѠ�F��>�Vv��<@�0y<�X�Ϧ�U+e��J�͖yF���2G5G�ׅ X�tT=��@����xA&��yO�4�Ԛ�R�:c�BZ$ǅ�Bx��/CN���*U)��s>K�(c\�\��9_i~�'c�+��pQ��u��� �s�q��gͤ��+���sPT�٨��񁰖�#�$!
��-J������{��z�Qݎ���}�1]�9�`�K{Y<��|�U�}n����Ro����դ9SuH��i�(㞉�|_������Aܐ�KK8l�����\pv��$֤ߧ�Y)!0�b,Q�)uO��$	y(��5��G(�=���D�V�H���
���ɀ_�0�ϴOFA@�';�������|��O˵����_�==K@-x�7��M:�\� ��8�&�\����l�|��e�=�����ޡ:,c9�ے��s���ht�����D����bk�u�t��<�e�Q�I��"�h$�G�勋��+�J8�
�C��V�����lޖ�{��e2<���W�����=�FOy54��fÿ!�s��C<��'���<��/ɥ�O�S���C9<8���@����!��]�"3�B�ִ.��y����T��f1�*�պaF�wҌ�h��Y��1���� #f}藼�ƛ��������xCb�n�ߒ�����!�ӈr�c3$��86f6=u�b4�ʃ��Q�G.�<O|�1:Y��!�ZO9�g�������������-�{�<��	C Ԅ�	�J��~�Lc��T5͠��v����pEQ�q��^Q��Bۤr"��_�����9��=x@�ʕ��ٵx��Υ�$ץN���/�,Kq(���}��:(��)�|�-�q�����ƄL��<����Wx	cd�a�|��dle�	p��a�NN��"Gd����S�2�rNl������6~�rêcf�@��f��(;��ƒ��ӆ=1OJ��;�r�e#<�A�c���cV�h��y�o�+���V�B�l9��Л*<C���~g_��A���2��pLҪw���,�������Z������R��?)������8$لQ;�R�M+N�M����e�0���HR���h.�~��S�r�V�nU��|��������9.�|}�Sc�J�|vh>�{F��;N;�����R*�����6ȃ����GAA68���Ӂ� ��s��l�86D�	��P���dw���Վ��Ǹ��\8��P-��is.Q4���:���%��gnȗ�{Z�x���(x��y�����pgk��������_��o�?���-��ݓ��Y֠^+�zf�ew�,/mHgqق���Y��4 sQX�YF��r��GA !��5��sT:���x���O��v�U���|JEZV´b��M4
8�۔��!��yM_3�x\\H�ۉ���y�'i��:)�g�k��{��G?���#9<�$˝w_�ѻ�T[6V5�����=
p8L�C��a9o���@�<ܴ���V'��\qf�Q�VΘKW�:%�����J��Dc�L. H�8`._�ʊ�W�|G��m�|WdA=�lkǀ���d<�����D#���L%�C�P�� �q��"��?�%8��*��נ�������׉����v����ÌP���g�契1'1�@@�ޣ�_.[;�L�ol�@"��������(�SQ�ۮ�z�7�yKt>�^t$vw)$w����ݽ�@���o�����0����m���1OɝF����M�m�̮_�Nς�%�܉����ƈ�R���p�-��]#6H�m��T�.,Y���4ci#������@1b;�� &�2sK��b���s���'܃�",�Q{�H���.���y-Q�;���E2��2Ƞ̙W�,��O�C1I���š2J��P���^��南sK�w-��AT�"�ȶ�v'v�A�Sb�K�9f���z�=ύ�#{!����9�)�����ʒ8����ҥ���0Ĝ���X��M;���-���n��!m�x�����(SQ9*��q%�7#�gr��t@����Z}<���A!��F�&�qZ�~v|z\jEy�D�Ԃ���h�+��lyb�˥�#�,�����[�G��<pq����ꨴ�<nc+Mr�3���l$��aniP~p�)����N�F.�C9�F��G��ևk��ԡ:�m0��c�u�'j?��d}yQ^��srv�+{����ƺ�j���� ��ޓ�7��ё���\��g<Ԡ��(S�uM����Ӳ���de�%���9a��ɢ���s���\L��(�&i�
�AT�H>���9*jX�4��p2B�,�	��ǂE/�O��������K����m��s�u��s��e�pvE��L������P���N������o��������}���r4���;/qr7�ݞ�J)��#Y^=c�Z�hǓ>yL�8	36�,4_c4"3(�R]/j��!J��'%���@�i��{�;�5��}�m�� �2ĜPك��ݻ���q��sum��'��fx��f{�-������0'�$�'#;�	U H[�zp�C����3���$4��������gT#R��m=��ߋ;:��@>~��Ju���������{0`����'w�7ei��N�&�����r���1���5�^��5��1X+]c��G�|��{Ӣ9�K��G�{�}:P�͸|�p��3�Ɲ�*�F,�{�����|1"�f�ET��zD]K�ˁ���L�޸S f�q��f:X㾜;sN�ٻ�,!��v�{�r��~N�D�f�:a]:	6
��:��cR/��վ���0�W�kR�[rL&��,,t�:��d&��6R�	dv]�cQ��:��%:R5� &��s"�"�b��F2�:pVds9�j)�z�/��8#@G�c�t����Z���Jb�:2��=5�qj����K<�^Q{��3�%�Ҁ����Iy��n�L�cL[�,���ѺF���=��N[�)x)����ey����o1:����Dƚ�����2���sR�yyדּRWf�4���!Zm��=�V�;��ZWh�&>ϻ'C�9N�N9�-gu�$
Q~QKkު �\�)�Մ:8VŒU�Ω���)s�S[K�0nZ���}���{8� �GCt�ޒ��)���7<��:��Q�����W���7t�)�>Mp���:89���ސkW/��ݷ�}$M��q�Iu��b������ޝ�U�x�my����-�B呞9w��NVp���(I^����ek��\��)�L��	S�ݶ�f>0t��_���������#���R?]z������Y�g��$��n�����L�d�ݙ��-�D�`=����W^x���x��-O�� ZYX�E�&��;������&�>qM���u�S��ߗ��ߦ��-�ѷM%��q��3D�.�Ã�i�fG����Knʒ��)�[@���@�L���4Ⱥ ����D{r*C��ZS<l6n#�\	K1n����y͐W�_�z�H#B8U�Nc ^^=f��n�3F��`C7M�{������[X\H5 ���0Ȝ@p�V�;�SDbf�=����\�`�{�Yb�H]����"f����RAVn���D��d=����,��8�L0=�f�Ƹ��S�f9�����s�2k0���N	8zXO[���>�]�c�{!��vj��T��9oS*�z�x.�~�i~����!���������~h΍:�V����Ӈz?mhH��i٠s��t�!���,_�������"whjT�W^g���_yMv��Occ�S�Ы~�|f�?�z�����?#ݰ�C����1��G�w�z�$�?:/z�@�� �S���kve�GG��g�������1j�_��_ʿ�?��%�a	)�4�4r�K�(#����/]�ٶ��Ze�i�De��b�C��ԇ��f�.(^����%�ruM�fm�8a�����������c.�կ|�+�|��a�͚$K�+1�K��gVU��U�]�/ �B� g4�g8c&�Mz�8ү�I��e��4Ɇ+8�`e�h�^k߫�*�-��������FV5�|h.,�ՙ�w�>���Ǐ�l�%F:�p����?����������+m�2�P����$��iy��*e��3a�k�������2)G������<yRN�:%��9~�8}��Ғ\�rE���ȍ��icG�B��ջ� ^��	6א�I��ޚ���(p�X[f"l����d�zg	v
F�D�\9�܃	5�b][s�� ?#���RO2��z� ���gr�3ُ��� �=ٖ��]yp�>}#�J�3#����6�m���[Z9!���*�>�>ς>d򓟨�hPa��Q�G�5jZ�UF
�{�	5�����7+RSc~W��>`-� �c��B��h/�O{|f@eh��^�OL<�H�e�2?La��88�ʹ� ���|�
P�Ҩ�A����_|F���濦=��n��:����vw�������ɹ3������y��������l�����QԜ�-���P`P��Wj!���������
�gc�3JU��X5���6oފ(��8gl\8,��f,@\]L0�[[y����"�w�Ց�.�0ޑ��>���lZ����B/�'� 놈22����b�\5R�zr�(�ܺ}��p#�z��s`Y�J\�u-�$� �5{��98��Q&آd�I����q��]�Շ���Uyc�k�XQ�ߓٹ6���{w�ӈ�����쌆.���yFE]ݱՍ�(��\ �k@[���\�pA.<�20��RU�&k�Z������u @�w���sA6 ����o��B�������[ ���e!�ꗩ�h��Y]�C]s��vF�����ə'�3w=�kx�ŗ8�	F����r����9Ө�n�e���?3>�#ϳ +֙c�ˏ>�] �H� ��.=]:�9���)��7d�C'뾴 `���'O�='������ŏ>d �	t�|)w��K,�+f�r�ZFŸ�����b��sU
����l�cv�֡w�Q{E�t�R{ϠD�G�<����D+�S�^:s�������[	G���������T�U~2�k������.~�1��0�g?����/Rw��}�����$o�	�~�?�����%N�>�S컯}�k� +�m��?��?�q|��?��r��V��V���K��o1���s�&BN��@gz�{�)'�64�J����Md7��jC�=a䇭<+9�
�jD�Bq���b�g{�����?�s�+��W�����DK��0̣��a�cy�`KԞ��@;Fto{GmĬ��\�rI�N�-RW_C��ؚa �^�!e��<��c-�#]�X�P��jƙg��)���S����f@e&�O�Ѩ�"Uo��k��ˇ+$=��ڐ��$d�b0Ӣ+Ks-�ҫ�#���?|]�
���U����ˇ~(�FS���/˙�g�3[�Ks2ߪIO���6Hܘ�����H����	]�U��D����wbE�{�Сb[�v�Ύ!<S��MLm�g�_a(�Ӧ�Q�j��΃�]��ݖ��%n���%^*y
��=��yleIz�G_�����K��!�+�+KdS$� �ZV�cu�����U����E�P��弦��i�GY�Ʈ��6�r��[���4��}Yaww;�����3����AZ��0�5�`��PT,f0<���k��)�T̜��AWn޸�2a��.�s�>��y*V�n* ��x�+��k�M9~F��
[���4 �0H��:�4���������bc>rz���E�f+~�8��H�n}_�TdV�a�$\���;�RK�ck�M�v�q4��=�H���,��Z���<���&�M���n[j��J��[��x`�	�]�����V�.����g�8�5�,u��G��w�$ZܤJ�?T�$C��JY���~$�������1����{��<�Q0�Pő���a��%b�7?�*�L8�JM#�����^Q��'_	�R��ڵ,-�Y9���gW˼�29��y\��Z:���#=�N ���g?�=�Y؂<��^Vh]�q�Vݹa}s�;���(_ xnHW�J�8?#�����VqM�;������U]#'	��9֗�,-k�+	tmR�/ƻ�~m�0h8C�D��?��i���׮�zo/����it�;q0��	t�����? �KґI�C�}��m�{��|�[ߐ��w?���}C҃�d���|��{ ���>4�$r��u�u�U� A�����OMT��J?X�ܳqʈN<5�{_�۸�ݗZ�z�C�X��HnW]�.��F���Ο9&�ϝ�˗.QEq8������,	�T�3��K�s�~��F����W4yocS�cCN[��̒d�Y� ʦ�Q���D�Uxx5x�ޞ�6�7��ذ	�up��4�L���#�!3 Z0nAZ(����7����������L��a�G��3$�~�7� /��"_����[o�%���ǉ"�U�C��;(Fa���*A����J��P���!�9[{*�]����������M�2�1Bh���91�� 1�Qq9�T&S��@�����u��TDG ����|uJC'�.�I�cf�P.��M�ҽ)�E�Gۑ�:d�&� @x��eo��Ӌkkk��Z�)m�l���Yw@�P�H�Pִ��E�	#t�E펕v��Z��F�6�Б�)~��!���6��$�>53�:��n(`k1{��9�<�j�y��'��֍�LJE�[�M�%x�`��%2���e���?�*�P���/F�ͦ֋=��`<A�Y��ՈʿF��A�s�r "���&tP^�ί�����6w�$U�3Fn�2�vfO�湢/r��3fT�k���bE��D��v������g���+�����lR�ӱ��"é �h$V���4����Ɠj�Ĝ��pDeW�B�+�̲Ϭ�h�8��4�����?	���txN�/1�!�����=��uϩ�{�c?;����됲G`��DL����(tz*�r̎+��@Z��M"	��Bܔ��C�N�?��=е����b��h��A\������ɉ����z=}}�m���0����,NS��cs5y��Y��H>���rp1w�ޤ��l{V���lo1cr�Ī,�,r��+ �޿+��ַ�=��l��T�@"G� ��7�,�:��g
�����9T�[�/)�Ju	����
��Ym����@����d�4��,5��$�:c*+��s����&�0ܜ?�7��.<�Tԇ￧AC�ԡ�?ܐK_�'�<''N��g�{^���9�d>l�5?&k[}E�#��J�Ya�%f5 }��3ؒ�Nkw��Rn�c'���yj��Q��(�p�g�%t��ؾ�:����)���ؤ[�@-s�|]��S�N����=|����,.��K/>+�{$�]�qK7�?�)�����C���80s�L��=҈>:K�S�٘�gy�ȇH!#���Y���gl|D�"����Ѯ%c����}v )@ֿң"s��4}Ġ��9re�Fd������&��5ΐH�2����������&�v�(f��}{�����~Ԉw�����R_|��<8�RY�����g��u pn,p����&��4ZM���U585ב=�d$����އ��h;q�&>��f� ��g�����!�ϯ�gT�A�z�XG�N���;�l���o^4�ZG"�O�ə�ڈ���6�k�k�[��	X�!3����,��ց�'8r�|�٠K*�����g���y��Ĩ�U��J!�섁�
����6m�w�Q �w���O<J��"������	��f��
;� 4�A@���ɂ܉S>!r��>3Z�%M��������U��T��j�@�26nX�$}�-�(�/�_u<�<���l��K�,����2L����2�����l������
<؅�k)�d�"�d62U���J�#D��0��GA�g^�~��(�>~�<� Y:uZ����:�s�z�	����:�1
���@>�}��Ǵ���~�)��'�Q���_|���dK�W_����O糠���d�^T���Ԕ�߻�Vfr��5RL�+�@D}
N�8�)ߣ�DI�d���e�Un�0���DçD7�G��r2d�*)�@؞lƙ�R�!����nOQ'ڐ�T�c.5�����մ^l���N03�鮡������uYԛ��f��j]NO��ș�����Y��^���3gOK�3������=l�5䴩�j ��ޒ�[�(o��}
�.��c��63+�s32P?��s�-��QD|}����v8�B��X���ٙ#D��Som>�w�~��V8��zο��ߐ��ߕ�w��6�reĳ�-���с7"��PCM�:�h�AO�D��U:�_|���;z�<�]H�`�F��ǥY=�쇿p��v�d�(����5��)�>}�O2herg�u�U�	����1C�@�eA��I]
Ό)o���j*����3��/��O�ΰV���<�j/<�RtT쾹�mt� �R���!�e/?�ڧ��ǒ�~���O_��!Sd���`w`B2]�zB��A�@���쇉�}}�UsnZl�}�r��W��usbNYv�'7ԁU92����g�>�fK�N���:�8�]��`D�B�����~e@l�HU�e�Nt
��dlS�!��t?�a�^��T}�$-q�D�M�H�G�K�<tv�Y�w(_���L��Ǖ5~��Ό��K1�~ׅ`�������fM4�k���>����<#}dYP�h��@6.bۮi	1��2=_�p�0�����D�7/,�I�VR�wac�Y//�p����Z~{�\z�k}w�o�.��p}���Z˽���F�s#�֡U�h: d�p$����A��L�1��y0����>'��>�v��
ٖ8�ܙ���o�,������K#Z��|�� �z{NFc謘~�����7k��۬���m�uG�~�&?y������?���9�u�lm?�8ʤ�ۓ���zj+�e5h��ڔw��!�r��E����ɵk��2�����Iv8�՜�me+J�7 {C`2Y����s��3�e�Z���~��Zo޽�f�� �29+Yu�5���S��J��u���w��7�sg�7^zZ�:{B.�;E��7^S�CެHo6!��6ww�33/�<��ܺ~��g�www_�V�h������P�]�&��3��:a�Mm�@8��.�~W�ѕ�
Tn���Hp��~��#"Imn^��F�[=�Y�	8EA����Ϭo��5�y��lS'��V���u^A����2
x{;[d�?�*��x�S}���+���c"t�t~�$���^����;8@�k!��z����}� ms�9y�'�s�{E�4|� �V1/��s��:O�3�X���u,����
�X����W���h�|�ӷ�9RcM9������#�+k�C~����v�s���ꍖM�U@�VV�v��y������97��_ L�f�Y7ﶮ�w������Oؒ^����.r
��h$}��\�|����.�U�Rd�ݒ�:%�ܼ��LTC}.v=ܸzQf��yz��(;���/,���WZD�3- ��=��NB�8�[*!�����gu����ٴN|	�t��gL�����4;�)K[y�!O�WFU���#7v^ߏ]C##����2s��՘EA$����ܴB"d�&0uޏ@��]l� Y�,6�%p����~�?���K�i@�F���֞����<y�	uL�,gvf��\g�u���~o��30[��H���Xwu^��M$'�[��J�$�¼4������������������>��h�t�r�$������5����gU�}A���ZL�����g2�A)�l5��J�t��=��'`���1.�(I����?��kJ�`1��J� �	+�� (���d8��[��!G��U)�~G2Q;�k�D_�vq�N��F��W�<>��}6��ܾ�������G,M�Gh����̲�z�ꇭ$8�O���59�z����g��G�.ɻ��X��۫sKj��y	��3Q�^Q�8	���t�`c����I��d�tѮ:+�i�.�&�!P������}�C6HZ�$CYX�a��M ��eݮ�s�>%�����|���9���S`��ŷ�8u�$7B���'tve��a��Z���~W<ܒ�̒�ӡ�����~��(���LA�^_c&pSl�b�W(���Y�|�}���`���nRL	3��u�F���:Q��袅3	ȒNH�2*���:}b��wF7�g=Z��g��+/�$��Y^Z��l?�����T+V{	��enF���\t���:�$һ�>J�Ӑ/~���sO���DԘʚ!���i�������>*� ���#�r��#-/��)���w��?�>V��(Pf�pBg�$,�����] u8��9��偮����lml��H1a�O=�2�'��� r���R�!��8hά?���/--��ا�G�,���9�Ԧ(uYا�������Q�4��a����s�p��7�>]�z�-�Ն�su<  j��.v�go�T&��Ui,m�:��ښ�#�Ǣb��I�"׆yx�/�o_�X�}Ij�F���˄���o��� 3Rb�'J�;]�rYЗ�L�#eى�Lh����y`�p�(�tX�O]9U��#�:�\τ-��޿�u��� '�م���BYd�F�=�`���[x���o��(9Q�(5p�N�/N�� ��sQ�940,�$�{���� ӡ��c+�x�L80�M�r�o0�[ϣ�����:#��ڑH��X�ྮx~�KBVǋ���L(�4�����θZ�(�9ˈA�Xj�����{E�8֚��R��f��!+�x �Pm胘���.�Z���ʥ�@�~�a=����P���Jd��5�a�� ��e�=���Xg�Cnmgt�̪�-�\ߠ�;���n���1<(������9�e{*����Җ@�  E-����	4l�I��f�ѝ��4�*�F-V2�y��䁯4
��byfV��ܼx[FM��a]._ o���ܼu�s��7�.p-���9�=t��+��ڪ; ��^�����Y=�;�=nH�6�=ߒ�ڠ�+bWc��궾Aݨ�eF��uPŜS�[~-��4�h@Y'�QO��J��>�Zs�n3�m����q���^ ��HZ�Q�I����{�l=\ׯ��(^�y�����Cy��ɪmY��ʛ�_��c�d��44�_/�qT�P���6���r!3�A+���������3\Zã�#E��&�ԙ�����{�ĩ'�Os�PM?wO#�EH��m����A�~���Tn$�7��[9;`k�Q��בQ���D�P��Ͽ,����
�θ�8�o~���|��E��/_�j�TJ�z~I9B*w��0���ŧc�]�(�xA8���PR�|\TN"�nz(s�k��ZzϜ>)����W ��~�g彏ߗ�������[w�wBghY���	ʾ�c:U���Bf��y�Xo\�&���l[�s�=����Fǥ�F�/~�K
T�������/꺾��F��r\�߿�����|�����َ�
�yf�$8�9+��5����۷�h �{��[k������9���hb-۩��ga�dˬ�3j��:)2���Y�Q��\&�:I�bsA�rĝ���ڃ<�S���G�-��5ԠD%]D�a�E���k�+;�)"���Q����⽑9#�	C�����){Zm�)G1�-����Y�k<j�H�l�32|��Mu
,;8�#��B�tz����$�3��y��➿;�w�>�Yޫ~?��B�:�
4>�8�[y��9gǑV���,�&�Fd?��׏�����CwG��kq��Ô�uR7})Hdp�R$�e{�/{�>�"��pl�i�j�nm�IO�I���yD�t��۰5��d�>pT1���2��ր�ɱ�u�'4��;�BzM��O������=�$����pG����.�j �V�sVP]}T���-���3����K����y6��޿��/��֎l����	�23��ΣD2�1sA\`�(����.ݾ�&{�C�{��kj7��Q�!�˧=>3������H'��3����vQr ՘� ��5���?TG�p`��<�-���3�rbU�D�=��������\$cE�M��)F���Pں��n�r�n�����=�ϜQ��R��ӗ�(�#j�9�R��ۑѶF=hS��\E��2[8a�
�"%���4SI��S���e(W��L�[�[d����R����Y��vW���$j*pkv�a1�4�ۺy�����M�ܳ��S1����{ y��̴]��
����ٳr���������84+��e QN��;ڻ}����r��g_G���*�W�3h�h�R��fK����=8�T���'Hz5���N�Ge�g�0�G�6�Ƶ�����:F&l2)9D����b'א+Y����w�sO���䷾�u���y���\��ʌ�~�6b��X�i��s|�G�5JK�h�\W{���F5'=�� G-"	3��=u�����;�`5CU'�F}�#Y.t�gZ<�ԏ�� �<<�-�j`�ʰhgG��\~3���a���
�Pxnԙ��\�d�rz�u��4R���ٕU^�9Pq��Mʠ��-0�z����Ag���?
�Ygń���=�$�=�ӥ3wn�e�I�ְm�-��HQn�R�Wb�_�I�_/f<y0	G@3N
�Iy?�M��Gs��ώ]>�~>��ǂ���Ӊq�e`�yU@����L^p������U�����9�w����C�ÃA�%St���ȕ��&|tyN�-�,��1C]�-�եS��fe�@&P�M,��÷���I��]�4� u9;gd��?��<�:����d��i`{��M}��]�nޑ�6�{����W>���o�)�VM��w)�u�����5a����%c��D��΢,��Z+$��&)M�i˖'�`}C�ܸ*G�n������?� }ȧ=>�ҏp��s'���x���-�^4ͤ�!�-���~��ܻ{�������m�K��j��V,$��G���n�tO�@S����>/3�~�oɇW�d���:����+���-jT�&Y:v�]6	tE$��Zl�3�Hr�iv�(�U��1�}@�;b�§��lA��ƭ'��,����ȹ�V�*�h�F��+�K|���w�;�p�nJ�ܬlnn��ڜBZ���y>z�H����Fb%0a�ʷ)zbyVO�<��qTG%*�m�=���Q������~U��8�&��MAH��j��f�ѠW\�i<����`E�%��GQ#��H5���������j�"Y����y�鉋��fa�p! 0*D���ϵ�7d��,A�� �HKs藥�9M|��� ��$B�,U�T�Շ
JV�*�Flo��>�OdWP&�д�;7��g悴�ؘ~�e�RtU�k�디2&~M�3'�k�sl \�ڔC�=26O0�`�'J���x`>���96�����|-y�{$;�_��}�	[Q�(��1��![:�Z
��w��a����@)}�9�#�-0:�h:���=����B�c�4`?� kƋ�����zғ��99~˟�e���9=�����{7�n-$2�or����)�������}������R2 ��
Y3?���9����Ey;5�!(l�?��o8��Z�6��i��"[rx��kn7mB72��H�䗆,{����x �_�dJ���{�T���,�;�.�'�4������L
F'�� �'�ފeF���3r��[�G�:��ڊ��v��jЃξ�Ƚ{w��ū�YV��{���\��#}�,_�dn��J�����D�����PD�pl��cdyKV`��fҨ�dT���lF��0�ɴ��%ȳ����t/L4��0�j�������e~�T��@+JD���(�WO�w��u��cvl��O�?��7e�XK>��Pn޾#�{����%]�s�;�g�Ѱc��ׇ^m���)"a�KGN*>�q�+��,'∖�M8���E{0�LG�C��� �o����/ˢ��ӫ�
~��{
�j&��7���|�6e׷w���(��[gÒ����n�����:	��E�A�2-� +\�H7�;�u���3&�T\_�)���mʾ����Pq���QB��r�^��ç�}����#�I�`p� s]PK�5Y�ȁ#{_��L�ޏ��?-���j���l�=0��.�ر(ى˗/��S�C�\�$�k΀�������oS��$吅i)����,a��@iX�9T/�=�� ����5B�!���G�\�qS���������<��W/S��	5�k�ڞ���N�k��9iɩK��Rz������QeA �ޢ��l�ŢtO����x��gV"���Z��"p�������_w��5����=��d���5���n�n�1�4��5��^Q%2��ά��.5�ו{����5]:�G9q����"[�����P3��z-��@�d "�J���`mA�ټ˗�r����C1��q>�����1�h%��Ԟ�6 {��p�&��C����Ϗ�_q�����o��k7�EEF{6���ky�y��e#ر�3�]�1߷��]K���#���^c�KlIH=�j��2�81y�f��~�I��/mY7��M��8YXI��'�g�o�v�VC~?�4�d��s�7�yƠ{����d~������=ɪ-��U�����7��o�L._�!�B�ug��� ��jC��@Ĕ�N���+����'$S߸�k�w&y�<����f� �d�誌���d��_��6u|vӓ?�`TO�"w?�#g"����ݚ��HqV���î���n�.'��FsF����s�ݸqKv��I�����d�hTɰ���B�>�В��}Y~������w���9�Ԫ�Y�h2Ӈ�,GLC(QD:F��)��e0�8�p�Dأ��k���-9zq�m����~�4U�[�8�9�w{���˿�����?^VO��V��9F�D'�W	�.]�*w�(��(�����3s����N��DR/%!3	�k��>V�&�9v���-�#���׫��Q�����%���I��R�O���ͪ���ϼ�����a�(I�;4D'����Bk�EZ7�&G�:�=N��M54��G��{�ۼ>d= Tp_�������B�jB=��#��Q�$�������SO�#C��>�z� ����񐚺if���T���d4���a������1�ʕk����F~�g���i���,��\����B�s['��&��F}YƃXs��}*G�&^�"�4���9���LG�DFl�� 	Q�)�ڐ�ݽm�˿�K�6}��yONS�k>ͲGη<��v퉤$�p➝<��Z�#�����b�Q�'4.AT�����O:���uc_D��,�@AAF�A�&��y�nA���.]���w�	�Kd hϜ9c:M����g\9��˲G�V���Q���e�����q���=���YV)��h��߿��f��,�W4,��U���ӗɷ+i�xm%�1}O��}���]�q�7Z^\�S����3�,�[�n�A�"5�
tF�L>eBo��kM�B��1�y�3�Cf�C������k��,�d�֖���[���*��]���K�g��_���%9P{u@ro��O{�=׶x+i����'嘾WE��a*���Q6��CgbS�S��Q�bg��!) -���<����*�P�?/Y�f4���z���Р�1�����i����:�
4�e���C����-y���am��33������D���:=>�fsVN�~BH*?��7H>�B��jP,��>�k,�%#֔�z��"X��iufڒ��� 4^F���3�U��#��,�I���4ޚ���9��;��������'I���_X�/�+�|_~��r����^��KgvA�zCz�;\��<Z����-���QNb5&��'��C�'� �{gj����oJ��fL��q�Q.�Xmx���{��-�(�V�����=iο�ڵ'9��;�ŋסm�0(�d��=R\���~4u��0̥�=���ڢ�̷�С��51�4Q�	�X.ۂ���_��_P���0n�w����rQA+�S��2H	�ޥV�ƾ�A؟�*8*�;�EmP����h��=����j�(k��G�G�x�b_�R�E���F�b��J6��1��Nd�ѬVYdj��Vj�T�<�I���t�	[�{tP�yF�`�I�=f����dT�HT��nn���"���wZ\\�ťE��A��~����B���p?-�l9�9������(�om
�>c�M���IfB~��)�8���ZܷKW�ȇA�AD��8��ʀ�<�K����}�	�n]N���{?+��}M��W���<��2��;a�G}6��{�#��s)}�Fq}�����݈�cr�`Oj��LGm�����{���ekc�NT d������1���P���$u��|/HQ��!��`�q8E��z������=�.�jeF���;+�A�b�N�<�K[mNwxY�F��0/� ����KA����,���I9�zN�W�HP��AZ��S��zOk�be ��/bP�ӏNI��q-6��[� �c��������|���MbE��#��0�p�!d�	��23�"{;�j���pcW7���Y{��K/ʪ�c�+��no��6t��;w��G^�����ևro}_��F�ۋ噗_�Z�-��RmuH�m�ZğP �Z�0�'a���L���Z�?�F̐�.r�G9K����k��@6a��{�$Ԍ��$ַ6�?}����}��e�����'�nߖ���3YS����K�Nh��`i��^Yy �Q+�Le�eF(����cS�ĳ�s���P�)�`h�46;��לq���?������X�M���:�#�N��=�F��l#w��<��n��ɻz.�َ�]�� �=ݺZ��E�̮N_�}�u��K��=����'���O�x��6���0!��V� w���y�,�a����+�U�Vf���s���X� �,	,�����Wj�����p�w4s�}jKDQ�ſ�����,"�e�
n���FiZ����?��}>�g|I���όK� �G���9���)6�\�ؚ���  �.�����1��K���xP��
fF��y�	 �U��(Ǐ�2r$(Q�ԫ2?;#s����h�"t�񕅥��%�#�9+��Y���tG�D��T=Uu#D)E/���)�U�o�A��.��8f^�\z�c�v6�3����sz+�^�Ύe���~9x9�����h4r �r�:LL�y�.>����s�}�ُRj��= @�������'!����n����=��a��ꛨ���0�v�.���T�>�h�O
���� ]m�5��^OF=!�d��KS�;��u��T�u�}��:Jܚ��:1��U����S��a�M񸏯]�^��>[<rd���@uV�I5�('����qY>���Ct�K��aK�Aw(���aS�,�z�!���.c���d�L���P�(��:pT^�{|1�]'�k]�H�H�GR��x�U[�6�~pS_�ԅ�ӍUQ���/>���~вYc:�N͏����@���GW�V���m�vj<z�,)*�[>A-�ꙌP�ǘ�.��A�-��o���`���02[h-Vx"��MӅ�H�"��Ɓ����R��j jX@]3P�	cuҋW.˕��d����r�:���ޮ��kF��؉Sj`Z��hd����mbf�̰sE���w��� ,�E�͉y�N#��@���*��n��GA�Ѳ���̵M���%��Y�gH\�Ń�tjNQt�L����w0��읎Myx$���l�r�4����P1�W6ޘa���Q����/麬r�r����|���!��.�7)K9��w@�˫��"�/_4	t>��r���o��k�P���6mꆇ{jg�#E��b�E`��3�?��D&R��ۙؼL}u*�����E".;��[�t�	�A1�8u��Y>����J��S��T�|���֕!콅%/<'<�j���SpJ�c}�������^(���o�$���B& u�$�RuDHyWt�=���������3�	t�-.�I�{���ڦ�>��@����5��C?�.��o/<w"ss��(c4�fńg�E�u��?@P8���-���k����:a�ȶ+����Ub�W�{��s�m���R�L}f#5l��E�Q	���G�AG������}f��1�G�	F�U�;AH�&�Ȣ(���~pY5dӭ��^�ZŎ���Ek�@?��4��h%Z�S���clSN�n����ɜX��qO��dwX��s:B�,Khvԏ-�0�����.3�l�ɇVE�cH- ����S/ɤ(qkQF�=r8*�UJN}M�Vdfn�]��X˴Duȵ��Sp�����%p�Ȟ�X@��Pv��q��b��DB�3ͨdA��T�e	)���bh�\�̓���㧞�C8غg:T��|0�'�M3�XN���S���g�����]�����k?��>�"Ac�J�3˧�ɧ_!:\��UTX�(; ���ҵpoHY�>r��C�-ci�/��^"�I|Ke%�f�&�5U��S���93?G�~�=���i{��n���	�4���Y���D���[z�sjD���M����1���%X���42�}L�"N�p����a�"wlH81,�ݝ���А%E��lL����Ҵ02>�Q��<��w��am]���k{dE��S7��~���9!�m�O���r��I^b]�=���O�n�8u8ם�m�pU����w��J�Ԩ� �E��|��F;�QZ�]��4a��-�;�R��33KN�4��u- MgY���A�'�J�)k���aD`��㹛�~�V&���C��鰩����/�㥔�� �����g0��0tJ�a%Νk./2ŧ�mG)+��F����l
v�8�LBf��VG�G0�ϡ��j�N�y�v��@d��Ad���ߧ�>�{�����Ͼ�-��z�I�}����3%6��+ǎ�4}29)3��(�������k{\Ѥ]�"��yC3Z���~�W@d$س�;�W� ��S
�,;��n�o�uss|Ⱥ��8�)g2K��,�y1�++��a�ѡJ��}�2`~Z�'×���I�|���4~��Y�TB+ybΤ?Qp�t��. )�m�Z_��V�=�{0	�E`[�, NA`��)8� ���Q�#`�w3V_i`,�A�J��(Ș�PR�¼��1��L*W�B!F����Ƚq�e� �}����7D)?�}f�9�]is�Dm�hy�@$�qxe�n���$��=�b�M�N��1����\�Z����8���$�\.AzK>�����X5�Y�oD�$˄�-z�|��"�mv���Os�<Tg�~��t�=n�F&�ݨ��#��C]p�_��N��N|�y��H1hIw?��瞗3^��Eu���N��=�,��BQa�kb�<�$���ɿO��26�u[d�Yy7��5��-��@�I��J��g�tf��N�ݬ��	P�BF��&���h��A�6s�M�x8{ �iT�Zm��0T,[Ү��l�E�"~����}:�텏�n�'�����*�Ȗ]-N�-'����/��n
�"j+R����Vż�
#0r��P�`M�����[5�z\���g��
��Qތ�-�׍'��amqbs����w)1sit)�3�*R��n<O��GV�����aQ�6�v䃏>fd�I�� $��7q��^�*��2m�0�"4 
b��}>�ǣe\�@dlY� �`����0\�vM����)��iG�D�k��<�>>;vG=�ٯ�r������V|���y�k�2�ͬ1B�V���Xm�?�8�N3�����J}��P"�ӱ�������C�g.<)�<���1��ƺ~�~d��?v|EΞR����{�M����I�o-�F����y��]F;Q�g���U���E�&�L��Dz�wx-�Ʒ��m��w�y�Y-\�ϊ=(���e�uU����,�21]�GKy���ye���G��]��J���`���o�F�R�eM7�2Q9�0����R\��Aw	���@6�����"@�� ��d벭A���
��XP�p��|G�M�]2P��cg�#�V 8����*2�+�~&���)��.�T��'1U�'�N�e�/�0 a#3�5�o-��@� �`�׀DC�vlmըKehG�h�1�`� 	U��r��.!�t��Ž4�z���E�G�8� *|v��ڧ���gTt���6{�\�$��K,լSW���
3
�Mtܜ>P� ����P&�r�aN�����y�;�{��m�'2%��}4V$<7��qY^���5�����=�xI����Fv��Ұ� 6����2��3�ȭ�PJ_�wp�#�g�.R���, �n0��6g7�@����PcR7/�b�к���=Xߡ�N���W�(�sѵP6",l ڣ���f#�Vp(��;d]?�ioo
XW��)����uF�����m����ӊ��].�$��k�F��ރ5��L��a\'O�R�!�/<��:�s������3*�s�υ�԰����sD4���|��h��� k���w���>���g����jr�)�2w����޻��Q=w�����WԦ�hpM���f���!��� "sH�2�M�%�3�N����y�8U���B���@��GR$�YI,���ꟓ�O⟿?r���,A�dS�ԯ߉�+��[���$j#��:�#��Eu��@�QӜ��?��G����Xr		��T;��� 3@�T9`�,���s��� 0o�Ky#���R���V^�0UӇ��)G֜��Ծ�5;GZ��Z\����ͯȭk�e��=�tr�����d.T�仠������I��>�m~��g2����?�\��O,�(��ܣaT���%����9 =t�6��G}��a�gv���<�dhe��y�L�Ə "_�)��-�� ��E�r�A`�%�,v�6�ٺј����qy��Y��cn��u���
�b4n�����ĺV1�C6ɛL(쇼PMB� xt�������k���|T���c$6��?U}�@f%'�D�i1�A����T�x��\ےR97�*	^k@�bLH�?�1*N�x�R�O����M�5��pTpi<�5�AA�th��a�~�4U��F��`ooߗ�we�!U7�@�I���@���ȴQ�-�[Y�'�~IN�}N*�Y���ARCZ����QT�,���Eẁ�\v��)Z��ד��F�eb��Rjy+�3�R�,>'��l�R��� "�Qh��f��@:�Ȍ?���3�MFpaV#���oK�,�����)h�m��u� j����~[�w6hdQ�I�:v�bk��T���j;"��M�F�#'�����q"�B�闔���,ĕKKyi-(y�2@�K�����E������7M�Jrh�F�y���҂W���L��:��W\�eN8�v�8 X�(bZ5�C�zV�wμ5?���:�`�����^��`6&�ٞ�A��Q��9M�MG?�,��f�*�FE�J�����H��u���H)������'�'$�Bbgg���D�y�:�T�}Ύ���֢�Mۮ�쇏�= �C's;P��4=�q�j�37�@5� ����G����B8��1) �٬�3�\`�7�]����٢��p���::H}�<�!��;��/3�\�1x��:%�lml�V`���=�IK�3xK��px�?�<��޸�ϼ�N����l��.��b�R�^�����c���.�c�?���ö�w��'�p�/��� ���9y*TxM���\GM~�H�U�t)z�~���h�>�y+�2�Vt2���(c7�������/;�����C�4�"��m���w��>2	|���(�T?���s>�f�g�	|�,t��2["���<q����P�ܺ�6s���-���Ȟ�dy�ekg�`b]�WG�jC2��g1���
�x�C�ͪ������du_�iG��d)s�r5��'�n!�/p�����9_U}I�2�z.��l�q�M}�P�S\����	� ��R��2��(oM�pa�W���čOM�=J?z�hN��c��SS�3��lz$�X05*lK����yi-,�±U��~�x[F�L!�M�G�_8{N�d�Oȉճ�r��`#�e�p������"n�>�`�i�p�W&w�Y��ϰOrPp�FK���i�y�ܓ�Ls�^_���c�������5�g�׃���l,9�����e���eE�[��+�BV-�	�p��I�3><L��Q��W.��G��6@�c˸`"+^��9�������xC��lo_&�5n��hT5��W)�9z�d�����$ruR��U��R暝 �i��[��TY^3M�΅�
��Ɉ��ea�^�*���s�6N�e��'_&��D��A.8��Rt)��RSv���炵��������tww���p�S�ݢCF���\[Ξ:!�/�/��=�~B��F���3P��YYY�h�E�����>dos����?���{2�߳q��0��K��jq����/푬�E��br����GK�̊_S���G1	���,c�v��4������6Ho{G��o���E���S�6��F۷�B��w����UC۝;w4�ߣ8�N�{ogǦu���>��:�I�	���M~�K?��O����o�7'�H�I��A��Qi �  ��IDATH��>���������,-/���˝[w�|������~�J���O��׿�+>S��cC��� xy�{�u�R���
�g�uV�)e�K= ����|�ߐ�^z��F++����?��ڶk\gt��b���J�Čb��$�걛H�� �(xh�z�Uro��=p� lG�!�y�;�\��~N��{wV���m�{#��Bj��W��A�m�Ci�<���}S��G��/ރ��8��T��Z��� r�׉�X�x�J�&d�B:G�C�2O '�$�$��O2G	��U*x�}}�Il��Z?��Yԟ����A�G��J��XX&4��%�jD�q	+t��M�`ς��E����,?.)�7j�]� w���<D/�fC���F���7�@f��kFÌ� D7�l�90�ʅG��	������F���Hj9I�]�l��n��	�L�A)��;dov�e��2$��FzF��/�d�0���u��������rR�ifn��L��" ��#�©�y[�ё�@G�	P���_�6��~�2I�Q4���Ǫ���\�;6�AvE)��n��FR o�<��qe���x��1��X@�yD�����\�Y�	)�)��8���H��h2I?A����z8�a@47?�����k78'��̐E2Vd�D<���}�y���o��,/�s& S�C_��O_�ݽr��
`���Uc��s��)�w�d�.˕���w�  @߿��Y*�?88�F��r�l���V*���D������{�L�־E�;�rIϯ�f<�֧�����>�A�	I�����dR���I�N�#!tM�̊���i��.L%d�E�$'wn �{ i�2*����1'I�g�U��<��4;�o�9[ӷ @�}��&� b��#�G��(/*�K������,�P}� 	�j�{�3ӒX�}i���(�#�³h/�'�o�	����`*k�2<vef�M��\��ϩ\J+gW�D>}}�5��~ܾ�����cJ2�7� ���1/K��uϣ��R(�\V2P�P//]����b����y�6z����p�0�{u�~��5�Sg��s �z.݉3�h�nXC61$R�6����'C��D�%�ۤO���١k��M��m��U�/�7�V!w���͆!"�Ԭ��:��Q`�4X�ku6
T���;�|/�)��5>D�F�"������?ӽ�4�-�'�E<�-�x�Oy|�@%J�j�&�v)<'�Dih�J���ґ�u��(Hp[Q4�q� $�[��]�uv )r] [�@���:
ԘO��6Z�4t�E2t�@�E#����nھ,��C]�/ml�+�0vx$kF-�0�YF1*S�{ �8U��p@�C�99Gq鋯�?��o���ɓ���._:Em����'�Ԁ��u�h��v���|]��'�z�[D8��=3(m���9�B�D922�N(�z��M�	�ᘪ)G��}�n��"p�:w��)�y�����꣯��\
�G�Ƌ-���cW���1��s�M�n������$0"��r1V{hi�̍�-�|�y$l���PC�)~�MF�<y��\�|�b{]pEEDb1�{+FPMMV��F�����_�'����?�/�+!'����Z�bݭ;�x�}owH=t��]̎"r@Б�=HP0������ �}5Ј�Вo|s��!�,�)���׉3���|�����ϑ)g������w��� �I�5��E~]Z7�$W����t��>#5o�"�� s��>�H������R�ס,z��%�?�o��57�W~���?�şˇ]��k�m�(�_j�ξ��)ŕ9��,���^��g.�l��aQ�c��P���׎�B�6#p�,����8Pb�CӴ�LuNx�p��|yq<��r�Vi�<���/��5��Z����5�6�K���%ә��q���w���⋖.�3�ߗϕYfJ�I��
-+��J�)��,Sƽ4�i��$���gt��+u��:����e8p/Q�Ō����,j@�\�w"k[r���Pi�m��Y` ?|���E�͢0[8��ȸ��N �$s �9�'��@8dr@�D��G��6�\0��T��q36��(FvM!al���n[z{�cc}�I_N����F~�:R/\O>����
���6
;.���(f�ܬ� ���eB�@#������F_kZzq{{��σ�WC�B� �"�F:P�\l5���fJ�b�z}5��P꺀:+s�>�09��h�"�E�3Hr�`ê���"6.
��0@T:����",��z�}��Q(WB������˅sgI�C4�4��Ҭ,��F�*�sm5]��"�7�ks��s\3z�Mm�ʎ(q�Yj�, b�����b ���΢0���hT2�,,2�́C5v�T�#\����=P*��9HP|&���1�\��k�fd���N� rE<���f�&�� ���c�URǓ�Q4I�ذ?b�퍙�dA"�ma����A:��F
����U��������T�\�x�<��Ӭ�_�z� ��@3��e1����Y�uoMnܸ'��U<��\��Cv a}�d�{-��ّ�Fl�S�98q̥���dqa�[�:��T����*xA�-��� <.t��Irqpn�L`Q�:Yh! ���kSY�����g�m�O��ֱ5j�!�ue�2xVj��@�?s|��A�f��	�x��:Fvľ�t��:C��֕�6������u�SY��:"L�����DbI�`�2�KҮe[.�3 y��mѮ��
0���oؼ�8,��,��g���dH��u?�ږ[w�qHe�ђ��)��=l�3��\Sd���/t;v����:6��W�{�5�A�����C��)�,̳���D�y<M���.ؠ���jNNwE
*@y�X��(e�>����$��| אq���(#GUdV��kJ�Y�� m!|Uj��3��:� ��ڌ.^�:Y*�*� C<7�n���e���siJ�3/��)�̪�C$��������>{ ��2��`���X�Mh��919I��,R���K�hb7O��0l���9�#I���'�s%�9,5��df<3ۃ�>��T�.2�K�"գT��Z2���Aow������w$��ԕ���8�U���sT�`}��mҊ��S'$5p�4~�R�t����y3�rh*8��!nllː��f��
0��x8bDp��+p� n8�Ka��.�3�(s���hĈ5�H�6ht���A��d�ZŲ0o���TlL
D.�NY��cM0�LmUt�V������y��Y:���-ޏ��D�gϞ�^x�_�d�����aݔ�gxݛ�];��,���[D����z�{.�١����)0�33FV_�H~��C��ڡ��m���uLO���.��q���r7�Ѵ�O��=Z�F�q
��7B�0�9���R:�G�T_ep@��� ��r(#�j�ª��)cD�s��Uu�]s'�<��������H���Y���8���A�<Le���*�����3��epQ�'tS��_x�%���4J���R����@�:M���\�u����<��g��dC�jq�P9�0��kZ"F� �3 T+P��i�N$�7e�@�1�������f��ҁwd�Z˙�l���$��m)97_��:(z��0�|p�ж�3��!խ������p (k''�b���g ����}`)�8�r=���a��h��Q�ao�AHʬ0�D~��]:�(A��ϔ�D/��3�$[��xMN�,q��tZ&r8�e7ۥ]�%�]��8���Е�
���r_:)��-e!��"���E�=_��L�I�e[�,�ѣL�-�'�������g���pB�]��Ȝ�dZ�&2i����w��5��	�|�6`���4��}��]o���Q#��;f@�ųG{r�%ֽ4u���v�?��	���DΧ���y�6j�P?88T0=8��#P	+a�ՄM&B'�Y�?�
��$p6�J���<!���-��$����2��{h�����.�{��SO g���
�ɔ��{��b|>��Q	��{�׆�2b[�Ԃ��:\�r��T�Ԙ6u�UÊ�AT��f��S�;V#�N�� 	y��X�h�Z�z�8��"�E"=��<��h�C?3�$�����ؕ�D���d<��,�;02�+�@G9K���w�xNB�֔��zJ�}�iYZ�WG�!��ߥSh�6Ý[�|�+_�����r��5�~�ll���:�K'>ꔜ�b֌�k�fù�\4�/�S`Ba([����_������dgg�E"F\�F'ߞ<��w��FĢ�iEY$����!�GĔ�W�g`my�d^#����hٓ�h��,1R�7
s��VP�H���g_:)�����>�� i�sqԱ/,/�gׯ�6.���Y� !�����k�t�����k����-��LR����}�[FA���(M�5�͍����M�r^�3��$Ŕl�ܦ��K�4�����z�t��5�ciap�s�b�k/�=X��N�<{V~��C:����+3�a�\̆As�	_������J���Gf����3�}8[h.�k�kR,�7�Ј�B�a�����y���0��2>!����-K@�%�j�EUZpa�(���Df�Mk�NM���ӝ�{fQ:�=��^Q��6t��2I��Cid�5C@���o�-� w8ʝ[~zP�sSص!��e��my�����Vu�'} R.�m��v�ƔKE�ڋ	�?�[��\�`��9Y�Wp@��R��OPF��2�-b�i�����>���m�v�l�����c�av<;���3Q�RM!-�!A7��y��`Yc���bI1'�H��iL GY��z�h� U����(]�A���<C�
)�1�4=��#7d|/d!����8L�h�b�I �����7T�V��3:p���0���l#8'�)8>S�2�`���%HQɬK�G��ی�޻��<L���a2�n�>�|R�l'L��L?N�0&��czݢ��LF�2�rbˏ� An�yP�di�z�}/Q\>�N3�XR�Hfi4#`%�u�s�����]�\�$w�6d��v����-���'�Ϟ��gO����W��S��w�uK��B�%���K�S�eƺwFn~~#~����K/$�RD���FE��:��<u@�l<��× �lO���߿r��U�G�.�i#u��ͯ�N�/`�i�$m< � ��0�o��&ۅ�&���F�0B�n��S`a���*(�T�����{�=���^����x���{����\�z��ۮ�$�)�]9J8�g�k�}�E&zo�}�v�,_��z󭷸�����`��������׿��{꜌P��(Aut<�������S�e� ��Џ�����l�M�N�#�lX��6W��$�e��������)~�>�o���Q�b��f����K�c�������@ �E�w"���W�~�e1ݝ�亷���h�f��"�'`�	�R���?��vd}s��;,�$Y�=��
|8#�@B�/꼜���ۂ'9�����c�Wk��I =���m"�x�áu��$l��1�K,R �<�h�s���ˊxnH9�u�Ov���IG۱�{����<��"^L�-���se��g�L� �؝[��	���2�5�q&��?�R$��=�E�����ⓧQ1	�H�b�]d�
^��s@k̤��^���K��|_7�Kw<�:N,H'�k�X\�r��a@X��-�I��e)�e�q�K�`A��Z�&�8\�0��]O*t|�`}�>ā�v����)B�ɭa��2���ً_��
�/֫3dU)�L��C�&��M�7�Lv~Y�:9�1Յ��9vc(F��(Z��`��:B|)�	#�d��po���q5vvV�柷@��]LY���?�Wx���ψ5qi����Y)����

������s(���L	�*I|M0d����	Y�����_�A����E���1v.«�����h�Ss�����e����O��s�RƲ��-7o���_����kr�:XJ��yT���^��Lj#0 /�����|���������J3Yν���>녅9*��/���O?M�ķPJ;�g���������A����u]dY$��\VЉ�B��5P ���-�._���+�?�n(`�П��ij��A5^_[��R��\�|Q>z�]� \��j��AD�12�)���kW��R�_�<x`���b�HCѨ�`�8<w�<ѧx}�"s�YL�t"�KE"6��Y�̔����{s���@e�7�~,����m���b�AH E�,6� 2o�����z���`tE��]kC���9U�7)�`L��^��]'W�QF��Ȯ�� �P��h8fD;�^L�dRf��tvDd�@$KuƸ�M�i�2��a@��2��8e�J��Eu��%~x_6�vy]x<�/ t�+�S0���&Y��S��S��Pa����S<�ȟSi�5��ۥƏdb�Y����e��~�3�{�7�3
�9i}��S�vӎ!����}XIS>S�fA�62�~V�*9��֬TZ�m�00�����P�Q0�Yf!gd4�w�Tt\S�I��E3q�J�k�e�2�(IEz�Xz	�� ��?����ʘx��`�زa`���0�*�A+Y4�S�\��� F\1��p��A���x2`Fg���k,"����� ��Z�q
��EAZϚ�6@%TGs�")�l�5���p!���,D= ���������� K�մ��xBr,N�Qz���r�;��)1a"V��D��#ħ��f���t2�7�������N��f]j+Os��@a�L���G�����X�=43T��N�����ׂ�n�I���esކ�H0.vd<�S�26����C��_�%7L��3H��I J.�������r���I�BGS�������L|��*�d}+��!�:�J�׹sg��z��d~qA����ЕۀL���V(
����w����,��AW�ʱc����9G�س3� sg��-���	p��>�陔���L��ݑ��8T��3�5jă�}%��� A�7CJ�K����cH�TK�Rz~_�0�����c�t����аxC��@���ܛ5ɖ^�a���+��[w�z��4 A�(�EKa���A/����a?x�����Y2%�"E�E� ���v��}��!3+�s����>��BC:�����[��y�7�o��^��h!P�<��x�(I�����^d��I�ǥ�^:��?g�#1!7�A0Ddc�^=m�/:f�N��>�]�Y7�"7�|q0�u���U��$���d���u4�|>����A��H�q����IN�X�O��X.a����GH?w�x�!�Wk��~�{� @}mlf��\�V�U�([`�]��l���/�<���V����uG��:&�������a|����ϻN�������"�����6f�/	!D`qN�j����:A�����2�v��H���\ 9Æ�%�ۺG��9z�A��ή舢`��^X-5���U��O�Ҧ��EØ��zH�-������Ƈ,Xa	ub�k��?��]�Q��NN �K�aߪ4�{F1�45NSb\��JRJ�y'���[��(Y�}����/�L� %�������X2�(�ٗ^eI��є�Q4�		󳴶l!��9�S�lnY
� ��W�}`��1f����0b%sP�C'L
h�U�#I�6�7��3)�*c#[n>�P�|�{��AK5V>�����]������3�KpL��{�H�xݮzDP�x�2�oo��|v떼��W����p�PjH��<�j��e�?�Cu�h�o���L�27��^�Ө�|�h��j\qN�^���{?>���>�����<��2SpS����p<s<���E0�%��V��7���ǟ�g}�"��������~�+_�����?��a�$WD&^}�k���O��G���1��FӲ?������!�j��%�{�=�{8tFz��jԊ$�.#��1R׃*�hJV��/7[4hY �YWݜ�;�?�j��jǩ����>F���Rfpt��j�Q"�����:��~:�2��LZ)==D�F��HQRF����q�P6��t  �)�����TI����x��m�`)���A�M���J`hq���4��Pu���"����z�iN���b�]� >��Z��$�gM�f���ʥ�;I�ʆ�73�~�2hΆr�"��l̩],#`���A�Q�>���sꄀ�dr�h��u�O�=d﯐v�=z��6'&f3}Ba�R$����dNr�~��S��45������M�Ϣz	���Qx�����J����1n�`��Zd� �T���:���}W=zp��,lx�e}��þa�[F�J�md�.C$�)RSm�i�~$�޲�!"-�s��RX/c�	)+U+L�M���8��X��PZ �C�w̪RT����MMjs��zvf�Pu���g^
�\�� ���6�N�e$�"�W�C�`�B�IЦ
{�b�p=���z}����sk�(�E���{\55����X1���BG���c�UQt;'s- �:}����#�ؚ��e�3��HL&Y' a^De�Y�. |.±����q����P�f:�I�����$�^}Ј�"*իwǃyh^���"+76�w��>��������r��]�������ŋ�)���[��Ç�I�k��;�?*� 	 4�򶞋ރ{�0.�m�&d%�����3��zOK���0*C��i�}����~c����+c"������]	��B܅ƜP�=�9#|�ϰ���#��PF�_�YX����S] .�O���Qv�	|"�݅�ez���/��?;��,�:��O�ژCddlE�ȁ�����r���Ԛ�%&E��e+�!��Z��`�P��?ֹ�`�4CD� ��������{��;w�����lA��xQ4*��#N���B!1���!x?��s�ˊ�3�)� W�Wp��#tq*R��l��x�����˵ ����w�=K������UO�K�f���1�$vQ� mf�s;��K'3]F��>e諤�=�Ҫ�ױڪ�t�n��3������%�~>��Q�+==@���4XA�S@S��h�U�у��\�
�wɁ���<��Q:��.����X�vp$�U�sl�~�u
�7���{�Q�,�|n�����Y�bN��;��;1Ǥk\ ��&\?�m��iO�a_�dݸq�<�S�������Ś��jv��	��}���M��u}*^R�v/8)5���t|p(#��ʒ��5�zu.2���N��J,G�#t(��Y��Y�^������VrV�U ��b����V�  �^�A_��tG}�y�X��H������(P�	T 0�8����Sgeu�-�I�ڑ��XA؞T[uB�[�JO����y`IL<� ><�I�D��C�ޭ$UE�mi��z}��Tz��4D)�偧��?;��t3P52��AH*	��V]��(�kѭ��	�t��z�}��L@n���'�5#M�
SLlW�o�!ԏ\$�I��@�	�H~�C�9K���8,��Y�"=����uP7��$iB\�ݼ-��ߗ_��_�^x�h��/U�|�	�
�x�y����Ͼ�y�����$��i�v�p��>{Jn`��M[y�$���?S�j���@��*R |�)9>VG�Q��a�8���"�郋J�AV�i�F� ���qw#��b��bi�q�N�7S:�������*���(�<I�|8GQEP�1�Z=�33�gVM]{0��jl��,ߨ������Q�$����b�OVF�==X�61[]X�7_M�E���#���\
��!��j=��I��@�Sor:�[l�$���U�i���ܿ'�����j���:�󝔂}E�}�imjz2����'�A�4�x��'@g�;��AMJ�(S	k�ݨ3%�D���=�c�w�2N؆�/���<Dh�wI�{f�ٿ�~�Z��XӸ�)9#�2�iJK�DG p5�C+��I��iW���bъU��V��%�  �T��is�!=�.$�<�Чc;��4���%��B(y]Aۡ����Y_�޻�*�L�i�u���I��)9"�E���P����˧!�W_�������7~���j��������l5 mA�R;��J .�|�����کv��i���c���riwl�_R%-�*��?'޶��Y�1�Ym�k�6�Z�xIG���3S��8 i��;ֹ/d��!��M*Y�A"�;H"(	�5�T! �ka�� XYhT������[��G���}�I��Y�M�DmJ�G��T��O�l=ڔ�'���!+z��'���׳�I��9-Y�"�8�S#��S�ʎH6�]+�f�� ��Y��짫}���U���iHs�l��{*!�d��N�N%i*(	�O}-�A�B&}�]��c�<x�@7_�@ŶN|OߕǊ�����;+d�/.�)�� ���GWf��!�To,0O�DE�9�)2=3�������J��3��t����saL�ܒ2!�#5V�M=�����;j�|�_�s<xp����ݗO?�!o����������{���*Kkjp��1�������T	u��B�1�>��X�7�>6� ��S#U�V'?��qD�E�
�o�>�������㪫8gW�L�Y��kAH��'�]<���`_)˚������2ea�k0�������;<{���/��z���F�z�*�Ѡy�?<�*�Ui���� g���mc�9w	�	����A���� R��CY)\��ͦ��@܄0�@���A|C���P�4͉j�A�K�o���mS�u��q�h�J9^��$?�@�L����/�d�A������9>�����6�Q96��q:�̼�oV>Se��6Ki��QF��E�r㨬A���s-YlUd}y^m΂,v�ҡ>�y� ���z(CF$s���%)�mB��-j&TŶ�Xd򣔨{��e�Ûփ�H���a��=\YY���@��o�AU����US ��Ęu�=��;�(MlcSΝ�g�i�&�1�}\��"ƣ/�{�>�ώ��x�O�#�T�Σz��^��I������沑bw HU �{��D�I�tݒμ��6h	�M���6VG���1:�M�1ҟ=�OI1 X��'��j{ED|�@V�$�U:�c�qcpNū&꜡b6�˭�?���}S�ޡ�l��� r���n�K҂�R�K�vy}Q�y��+X��ߑ�n,����"��{����=��[m�����$�WX�s� J�he�\5pTM���&����/��y=K�A�EQ �`p(p���F�3�G̹�Fq�ޒN\W�ޗ��n�K�=#���_����_����Tm5����rm+�q�����e���;" �������O�JF��$�Ł�8P�h��y�d�KٽB ɞ���^y��x4&��<��.�V�ҿx�uy����a�u;��>����{��`B�HN)��8�g���\w�$���@��C�G����R��6o(#���p�!)	i���5{��!S�1n�� �����.��'��@)U����ɞ�ς��K����V��΂�Q7q���H;+�0�1�l�)��1�o��R�y�F.�z�)�q`��C��Z�B�� @9+��4�tNz]�莬J�ȿ�{j8�ǌ��u:䨠t��5
D����8H���
3'֖�=}@�y�,%� R���l�u�\��M:�y.�CҤ 9�s2P(�P�0�A���A��V��N��|h*����Rl����������;0�7�1�f��[D��j�Y^T8,��b|T�&�MIL�v^z��	��ƨ��&�"<�zP�����& ��ʘƃ�٤RDO�}$a?�ۢ�����N�qa�!jO;g�z�u��?桨p��7iU�-*��78��ǌ�����Zvpo֬� A�����C��-�2��0Ҋ�D�M?/R{���{Lf���o���\V�E	:Vs���@.���fֈ�ؐ���x$
�)p�x��M���lG��`¶
��Z���D�pXO3k��������WM�(� �e
�&��D����~�p�c\Þ��H�;�G���{o���^��:��M]ǲ����:�N��l�����i��v7�ʙs����IcqM��Goˤr�g�Ei6Zr���+����Z0h��a���d!�����gcn��??���|KG:�	��fܹf·��F{k#ݘY���2�l �������\��!�WA����Y^YU�f�ߑw1|�#=��F�{����eY�_T�v^���V�Re�g2�1gQ�9(�I���� ��Ag	��x�̳�!�_	��Fd6l�@��Jl�3f��P6*,}�W㵵�-=�fx���0��f(Z�|���q����Y�[4/&O%t�1[���Xl���!
Ð����!��M������v��F*J��4oǉ���a��;�!���^�����a�C�4�a���c��̛2g�Q���{�S��S;D�d�,Ȍ7���u�� bq��,�U��Q����{A�]�sT��h�'=�Ի
O�1:��!�������X
J?�P�~�c�������1���A�ظ/�j�?	�Pƕ��-m1�an���V\tv�� ��=c�I����<��Z5��2d�h|�*��ߊ�E\ Y���ԋ��b��p�!Æ�nmm1}�+�7n)�I���a�������h��?f�tr���-)��;K�<��HԱ�.F]?�0� � �� � ��S�h���tR�-�oU��a+�$�	�r�]y�B�G#��c�Ef)�z]=X�.��kMFS����'9b�clh�D@���\m�H�VN���ȣB�s���~y�9xy��r2r���u�?w@���Lº���I`��Ig<���RT�AJ�"+�7±$���v 5D
X��O��kmuU��~��UW�1�ձ��1D�b1>��X5D��R��FϾF�ML9=̲���&�e\c0
_ú�l���d�=���/��l~���<��}ߡ�0�=�{++�t�!&���(��x��m�I5�s^�����փ;r���·�r�����������Á�FВ!A?7�fZ-%���k)�����_��dN*Iq3�i���J�U����L��H�����������gפS�o~�o��w�#��1��ȵw_�y=�R�G�PP�`����hoK͆\��=���jUm��>&�0Ϫ$(Q����W�ff�gb����(b�1��8pf��Yo,<ob��ظ��i[XZbx�,&�"GZ#o�A��5@vSn�}���A��j�P���z3���=�Q��9*�麼��G�W�,+�1r��̉��F���m�?_�͛�!T�Q���2�E�xJ��3܏�J���I`Ŀg����4�9��R7K�c�qC��q��P���1�댪�9���
: ��C2 ѕ @6�
 0V/��s�V�_�QA�����S-D�J��3�A?ßi��z��x���h�6�\��+NQގ��$	���u�x>��ʎ�i�#��1㹺!矡��πF�hQ�/��x�x.�6�>�X8Xq���[*�p�AO�Hz݌'Ђ^(5`�p�A�
�$�"k��*eږ��z��#�����3�w�s���ba�F~B�b@��W`
e�Ct G�xb�S��/"D���}��a����TA="4c����!���$G��_�#�|4��:a�R�I��7�i�~]��3g�竄(-9>&�EP7�Q$���G�h�Z)���9L|]R����]���P��w M��4LE��&#�V]�s�I��T�!jp=��geqAV�`�*,���o�u@W{�QG���G��<��5uD���:����,%PeO@��gI��W0�$��#;�u_��]�|�N)�x��5ټwKV�;ҩL��S���Oʯ��e����viog�ʙs����y��������i]�����t�6���%o��YX]��Μ��t��fS�:��i�h$t��'��VVmq}� ��/�D���Υ��˓�Tp���}�,�|�PZ���Xr4���{7��wߒioSjKM�lɸ�]5o)��_�W�G�6w���[r��tգ��?��0��|C������\}�9wzY�o�$6�Bf�T� )��`�-d����J�+l%��S�8��a�3�K?�����"K�lOB&j5����7fth��2��q)q͚xS)�RR�{T�(\H�65�fx�qgjޑXQTS�r�����{��d8/�Л�g�{)��7���H�F�G����AC�Y�R\�:*����[�̓*i����x(K����a�<��4J��*k 4ү*�ƺ�6t=�‵m����(��uT��E���>�!7�_�C�#�IB�oso�k֪Ȫ�^^�anDA��fAqj�!h��t�������H>�C?�c�R
ǣaa<Qu��fDgK`��E���G����y��P|�8~(9���Ǉk%3] k 3̋�d3�������J�b�=�h�o0p��
�F荥c��P�QW����̃����|HT$Vj������4�����+-z�':; ��5EB�⥫:ދzX���/�!Ғ���vyYOР�]����}=\ NY1�����k���կ~U��?�'�8�]Q�م��J�ݝ��#>g�C�sY�<D6�Xs�F�� JcN���$/)��PsvpT��1>�OC�v��� �v���&�Z�}��S؄ӄ/���/��5Ϗ���da��S�r�c�����w�Y��W#�jO�$h�5��LY�cJ�A����iX�>Ţ���"k+<�-)��-�O��箞����p��������ԴM���`Dpu��$ڛ��+��Ïo�hؓ�Jr��ۏ�ۯ�H���B��ã.1I5]���eU�pLٚ�D$ȁ��=��7%$D/���'�O&�A�˜���a�X���F�`*߹�������SY��~�}9�ږ�������}n��~u���~��E[��U�aB���ʲ<|�+�~,�g���N���|�t���	����M�H�ײ{ڪx��0���f�n���Y�Q�Ѐ�M��h�MG�h�aA�ܧ4��ev;���]^�����k���F�����U^�U��U;�g��AV���ݭ�pP�lnnɝ������pp�$<�J}6��cϹ{\��C�Y휰���O9��5b��B�A=U�lv�f@CH���J������|�ފ?YI��994��8�!�~8v!ՂJ�J�S��%���܀�`�KܨSr�s� 6�i�gC;����>�G����s2P �������� y���Q^�]2E٢����s�Mp#ԣ��d��Έ�4�n	矸�{�3��[�0�x\z��}<{���=c'):�)����4�*ѩ��y,N��,t�������9*������}b����1�w�Ѧ�.���:� �����m�����BX� &!�������¼\�x^���L;{D��*}��AO��r�{�H���r�U�Ҹq9��2;��=����+JXu���W�K_zQz{<�0�(��&m���ָ�j;��0���������������Df�Ss�zJ9
�{��c�Φ�b�W�t�Ƕp��63߇�;zM|�@?�s8H��f��pP�3V�I)|�� ?mPdt�`o�F�w�h�4����Z!AvjoϞ=�(��޾�m�s?߾��>�#!i�Ϝ�Y,jb�
��4�0Ɨ�m�8���)��.��A!����粞w�:�7>|O�����ȕ�EYlTeI���b�.{~�MP��>n J,YV��^�+�/+8�dKϚͭ��3O���H����r��g��ދ�r�<����@˞������,IFy�gA]>�k�Y�$D��1?;N��{���Lt��p���%�~pc�$w�s���|��;��Y�S��þ��.ˍ�>�G�3_�эO䓏>������{@M�#)��4�:1m�s�W_~J:��������Kg����+Mhi�GP��
��EY�Ԙ�Aↇ?�̌=m���B�e�T��
��8�Q=��,�L��px�.-ˤ3�$��{z>X�+ꥁ��+��TCר)�������2��]&�������!�ͺ����"�@�	���(
?:�*����LH�qV
���q$�s ��+���Ů\꩝�#�ņ�)³n��`���u�!����Cy�����R7.ƙ3���_�ȞyŪ���#�R-9��23
�%	�,5��|�ҩu��AbR�+��	��@���1Ϙ���{�Sk����>����o��GPR�9��{�;��ߕ���G���(�>A�B	��rK�e-��:��#�L�$�͵�\#���9s�����߰,}��ݻ'ׯ"�~��:
wewoO�|?��<\�n��#�������0���#�Q\v��Q/���f���{������~ b�V�����8ϧ��'X_����w~��T�'&����+ۺ6ۋ� ��gS�q���rj+W.��z ��$y�.k�O���r��A���&<�Ȗ�i؊���H�QPe�d&tA�7�+��i�8X)8�[��"0{p�g
HItZ���qB��P���ʥK��YQ��1z�7�ߗn�:3���GF� @�,�~o!}�%A�˒JE���8��I����f٠��W�)��t�~�)n<�v��[__W q�@���ݿ�ԇG�(TG.O]�un�A���C�5��"JЃ��cK�^:���O?�D�M+`����A8K���Bvz��G�k��9I�kX5^P�ł�Pg���n���.�4��TZj�V��2�F���@��ŗ啧����=���5[\��V֒�5T��U������(��F._�*�;{r��G���+/��
U᧓�\�p��)Җ�ߕ�g/�miS�`4>ֽ�v�����Z��-p�ơ:p*��L�����ד��稨ϰQx�u�*�j��!9�g#����ɝ��h��	bu��y#`���?�c=vu����ot�m�ubգA���Kg�q��hɷ~�YYV�����t����i���e��p�CYk����2�>�1��-4=	�
%zݘ��m��˯X8,cYYf�'֩ղ&�z���96B�2�n���=lRi꘵���Ѷ�+�K+D� ��&��_GT ��'�	�����0 �܂`Q5T98��SF�4|��z�v�����ᣇ|�$���T��y������њ�g������u�1�����x=t\�,��W%2o.%/�d����Tu�b�����O�TQ�}ݸ}+����؞�F�.�?LLD��,T��.����yXP�m���~B���}�p��� 0.󪰉S�ҍ�t�f��yF�r5�|���~�@�����{O��+�*{
n޽c�t(�&����D���O?�F�@F��x��{!�Vg�I�3j؟�9��/~�z1h/�ʗ^�?�.�����-����J���MIvGEP�V�A�U�l�>g�R1���W�>�م�hG"}  Z��&�������@^�޳k|�J�1=U�,/.�QUΞ���?��d����w���B�R�(�S׬���azݪ\�y��T٠�$�1��0���SmH1��N�z_=�d'��,� ?����	K듊�	5u��*�I�	JC���`�h�.�쒝�~��7����9�!���~M����[�y�5v��}�n�>q�J�  C��k��_�6]�R>!��2�_rü���)_��?����o�ڜ[���⨊ې��|?��&����(�@˃(�yG�B����k�X�F��	�*���{Q�W8����l߄)�s
�Ǻn��<���{��A�Ov 
�� {;�� ��Lx�T�1�#�����2�?١�ڒ��W�������z@5��BSGn(�V*7n>����'�\T�Z��w�A���S�pܿ�����~G���n.��;��꼧��:"���U�x鲼�ֻ��MYRp������]9���h(�jT�����H��8/YZ:�<[*���&���T$�|�?_(P���Y2���Ό�9�!eU��N�Pv�e��tv�^Ș9��vC.\8'Ͽ�"	����Z?�M���RZmE�����Y_[�'��4�yt���>~B�����7ޕO�kܸ���|���^�#�9q�2��xE�s�=vi�$�=��"0t�rA�P�y�'Ȥ(�MCKheLN���(��9HM��@hz��^Ξ����"W�^�-� ��?����e���܋�6ù��3Q�������Bw�(=S�����)ڦE:	���իO���L��J�+�t���ɬQ�g�ÿ'I�qx�=�8��i)P�&6O���a�W��#�G�cB�f����Prk�5<�����!E��|M��'D��{XE��k==�dZ3�\��������?�X��e!Z�
ns��v����)��y���8ͯ�����*e�:����կ}S:�Ի���� ǜ�������:����AQ��y��Ctǁ�5�	�^��N�S�P6��P�Hїk,��R�9��%&M`5/=t��2�W1A(�Y΍�T��;ǩK_3��ar���
��0�~J����"\-�<%�XҹVOM�~�Y�J��S	` �7J����G�"*�D�/cϡ ��H�{���5��%���g���k���Y6�ƪ�g�A!��U
�C�0�u�� O�88=m,uG}]?�_\O=�,	�L=�}om��wzLǱK���E�d�T-�Sڼ(}VD��P^��3_%�.�I�`'&���ֈ�������5]�$sg�>S�,�����\FF[�@@ ���}*��|�9
2l�-L{�4'h�$�F7�tR5^	�5ټ{C�n}$?��{$}�i�`j�����ūr�ѐ�)��0L�^�]��P���DAW����l�d
h��=���&�p��,,-��ϔ���[���,�/?)��k�F9�l2�S�jV�1F�}N8E���:J=jU���Y<W%+��Yt��[�@{=.���/:��N���ߨ-���(��������f���-̩������˲��!J��!�PH�k(>gog�y��iy�K�*�v�<��W��_�O��{�����øYSk�TՅ���0���A��a��7���8OC�@�5�̿v^�	��ҌIC�,-v䛿�zxˋ�/뿿�4&�܅�2�G�����ǌ,W�4�lf�\{V�����a�����T���r��B{;�]��yj�l��0�=��ͱ�9*��.��ߏ�.7�'��sT&Aʺ 7H�w{V�����*��$�G�Ex���z�Q�#f���fȃ�*�Ǉ���X��O��<�X}�*
=��6eI��i�T��1���?�͍5�g�hS;����余<D�V�}�KE_x�yV��bn|^��!���5ż=�+'�U��Y���EN��`�P�$c�ʌ9�Fk���|pm��;
}x�����#D��U��o��@�e iZr0<��#?���}-���I����GqQ�T�)p`����/J��d�Ee��^��׬�oT��y!�7�`hK�<au��)4Lz
���GЈcb'{�`�p��ƅ`_8	e"�4Q��'�����T#"���;4�`A�;4ք�����>כ�T �q�Y'c6�b��*&�~�r��'U�����G�Tx���x�b�:�������qŠ�m|Y�V�_B$��ڪ�;��S_��۷����Sʰ��6K�����Y�v��L3��}͜�[��e��u^�,�\�4mnݔ��I���������IB��O��kuDp��K��#�,�27>����P:j�V7N˾��*t]��
�� �]��=��c6�<��u��Y��I���X$�|aR���D��G�?��/P �$�Vy���u4�#V`���M\�9ߜc>uU�	6���2�0� ����{���G�y�v��HJW�"�"}zSzê,m\e�ﾢ�S������:-Qb>����}�}|WƃC���MsaIV�u�����M�T�����E�d�i�gF�:4#��:� �>�S>�Ǐ�҅x��g�0�V�;/���wdG=����#o}p�=C���'��͒R��AJ�K�^� l��!�Z��wB$���� ���t��<��?����I�+&����s �F/%���Fyh!Z��wr(�
E�R�bTA7ރ2� f��=ҩs#��9R\$�NG��{ɢi�a�ȱ��� �zEs�i0~h\���ޕ�?��<d�w�pt�mnJka��m�~��'r��n�ʯ~�)�^S�����s��>�}0��t�����q�#c�cc�y=���T�h\��Ɨ�c�A�n��id�QB�x�)����q��U����Y!�N~R���#�Ȁo㇣�G{DI,m����*��а�@+Ռ�;� X�F�칂S�D�b}�L�*��8\u��w@2D��;��\Xtr�G0��X�6�^� �iR��ZJn�<����oFM1Q2�m�|]��a7u�M�\����x`$g���,����\NV�p�a�c�/�^@	3�(y*y�A.���Џ	���8	���؎�'���;���k�݃#�t\�,�c��y!b�}�%��>�+����u4<|Lj���`p$9�Y�	�1�ء�
�\ޜp~�g"u.���gNO��f��v��Lg�%��lCn�p^%1���=�6Նq���O�Z�W_~Z�=<T��啯|YΝ�"���M=/iS�7��{��`�';ۛ<�����q��e2�'ݣ�Ӻn Ъ����k<Z�4Y�OJ�_���Ym �s|�n[?;Q�*imX�U��J��)���+{�ԚU�c�7� ��Hj��Ԛr��ey������_�����3��W^�y��Y�*��l�<�w�}Wn��D=��r�ʓ�F�m�XW�)�F�"C�N ����=�&H�m�Ӆ�C\X&��F�u������o�Hz�'����K�Lv�H3�?��^��1`aWVV�1�sL���x�d��a�?ȃ�|��@���n"��ƍ�ab�P��nD*5C��P�����[�^+��ٳ��K_z�<��߻���I�'.<y���;���W֏�Qc�l~����Bp�&d]���o�XX����K� ��*�l4�N��M���εζ'/+�Ņ�B�@�����SzY��z �Ω�USo�C�6)Eذ�'��L�v�ܻu�@H�o>zȦ�&DϘ�>���RW��l���}���������{�x��ӫ4� .�Dg� %�����l]�<50�?�xrd�Ԝ�u�ߙ�
)�l-TWMg7b^=�T+��_W�9( �^�
C�H��TZ��F� G*&N#�F<��J�z�
�ź.H�&·�T�3�a!R65�Q�RK?�� @�$&��qV��"���`�?K<ʒ���$�\'�=z,����+�-Vk�I�O&Vjm^o�!�B4�xo�I�I�n���)�����$�գ'�O�W���ٽ*'��)���S��"��ː?/Z��~<~q� ���ؙ~��{[J<3ݢɄ���ɖ}rY���ql�c����{�X� ��-a[�I�ƺ��s1�^C��]E���c8�G��v|@>�����N뵌U6����jIK��!���l��������oU�o���_~�2�KkgDc��F
�P�WS�f���9m�_�q�jaM_3"��+Ic���y��ĜM#�}��[J3�y��K��J$��7^䚁��pBQ�`��aU7~��Cx�+�kr��C��[<}f��9x�KK+r��%2��|�MzXcE� �>z�?_^ ��Ey�7*��Y�8�<!j4@��~tW�+H9>�L�&�{r��֘�����IY�w24�o�Ƙ�k(��D�������v�lȕKB^��͛&D����'������<��'���CьO�Y�ڨr[5m,V�fia��t�4K���������z[^��:�5;�C_\'A�D��8�_'��_�b��@��SB���J/ID�>Sm�K6Iua�&���q����d��-,B�CR�����Ӥ��d񐡑^R���1� �����;҃���ˀ��u�Z��&���ļ�JMe�sV�����?���G<h!�����bF��Z�<*��r���]��:Қ��++k������@a�B�$�*x,�a���p�q>B�Nv����X� m���C����<��89��gE�∌�[����u��2Ƅ�{�L�m�W���,MM��Wn��D{���Q���Q��-�ϰ�A ���z ����|F�
H;���?<-�B�XD�B�\��|�%v��h,�tOP�vJi �)��\3ED�ie����i��R�t�V��>N�4(Z��G5�=��a�.�k����~V��L�|��iiO��=ǽ���6���1�*��Թ��`���`od,��Dxa����Gɧ�~&]u젥��8X����z����ϔ���:��`�t�q�X$�,�Y_�`�Qߑ��Ȧ�d���B�@�������ẍٛo���禼��۲�w ��EF<P�S_]���?� �I0`���$��เ�z&�b_��Z��z&V�V�)gl�����_J���Ǧ�b%�G�LZ;�����iX�5�PY!Rr@�̍;�s��d>ڔ���r��W�ھy�3y��r<Jek���'���b�h����o~]�:��_�/;{]��9�)�n7,j+�h������Lof�1K{4,%��@�Kg#)�b��^�I�M7Ȑ8��Cv�\P���	���z��(@��;����JNx7I	`��ȝ� ��ρ�?}洼��󲱱���)�@�V�
�}Eo
�M˲ē ��7�wsr|�Jb�u�Hѽ.���<�Nm��K��R[��Z|*�ppudq� ���)Y=�ο����Wރ�s%��C��"J4����<�`��Ņe�c�U������G3�Wa��<I���z����R��<��N���
��ҥK$ā$�vz�����:a%��K�&˵�?нc<����v�(")H+�aW���UO��<��+NݔJ���U|ZpD\,���$䐨�F��8��D �%��R��9�M�1���r�ĵ�g�e�! @v3O�з��Rao*!z��C�cx�*i�����I;$V	6a_�[CP\����4	}�0f�B�d��J�߷x�$$���ȭ���bd�L���2#է�� -�77�����}F[��0
-p��	'���?��s�'�YL�Ņ����aqN��e��+���sTf����S_3�,���Ec��j5�����Z",�����9VMK�H�?�]�߻�G���љ'Q������3��>�$�b�V�9_9m�q�ёL�5�N]���ҿv�;�_�CEG���	� %�ߑ�n�}lu�w8�[{j{�k���G���v��=~f���g䒴h�"�Ρ�>%����Nm虳*��~��xH�xQ�N��d�jϕ罞DѨ8�E�9��%Z�0o8!y�/G�'�7�d�e]09���ʱ	����W���R�@
CS7�Z�_:����4��l�h$osq"��/ȇ��,ȋ/� ���o�{�?�n�ݻ[$�U͢�f=+�Մe�\����g�b�S�nFl4�����I�3+s-	e�H��R��FgW��0��� �T����F�j��%?.ߛ/a�H *fh�J�2�mgW�SO=)���}���^�߻�@^|�%y�h���_c��I5�)>���#�䬸�3�1�����4�)J8�G��c�J!����/��1}�����W_������Q�����K�h��`�*�IOn&Ĭ��R0�N�hH�����h,�R����}��Ϗ^��u�5q��ت5��a��9��矗N��T	�} �Z��
#9�[���7BɪU J�c��@4_^��~ʦE�����g&@8��|U������3���D�	��b��h�޶�������LRV�
��x���������x�9��u�"�2%L��Z?ʹ�a����yH��\ǥ�� 2��㐁!H�Vr6)\ҵ&k��:�Nvu��'J�'Y�g�
ʓ��i�v���</��YRYM�=��&솋(	�n1w���MVM]a4�������J$N�Dz(y�L�cNZ^�_bN��"';�{z0V����b!>_/�NF��z?/{�`�Oګ�~�ez��:��L	�׼:�G2��7>#G˄�+�ğMFSs�Az��$��*�kT�DYLJ	DZ];s�y�W�p��Ŵ0R��k��U��]܃qI�e�=ϵ�W@��s$���������H�O�M0sQ���{�߷��gO+`i��;�!ѓKW��7������-�q��R���o�foo�0tbϹ�s�lP�����N�����M�em�nȜ��J ����!jH��'��!��uR���7v���d(�U�z��u����=VCtǁ,�0D5Կ���ݶjj�h��ڹ�-�~vGv��R�os�-����L��������	L��>��'R ��%v���̿�S֫��45)n�Y���(�I~(���<9�~M��|$��ߵP�~��WH�:8�RNߍ;=Vz��Is�Y�/��[�B���s���1\�C�8��K��\T�����nm��wC>���
5�P�C@���k�#L����P'	�n��<�wc��'柍�p	�=1�y�|al�~�Iz ��@�
�<Gc���h��B�j���]�T&��UB���A�	)H b���������3�5ʽ�Y��$ ���]���}<��
�!x��m���MaW�
<��+B�< �����8K��2�Zi�dq��7���?T� 
i/둖+}d%� ��u����6�<)e���&�7?ocyL�|�u�r�,�&�e�j,����$�ǡ^x�~0[�#�!L�p�cD���S���/<G�i�g�~X+G5S7'O��*��c_�|�g2]�w�dA������;ʽ�Y��;���[�`k[�pK�� ֬�.��O�5�>a�n��aSZ�R!��R�5����`g�{]�Aޕ�u��Ҝ>��+�Ç.Ӟ~�h�E��,�����(��8�R���t�������	��󈩷��C�0�"*��H�ȹm�?l]�FCV��T��� �
��I�yTM���I$X�Mm���D痽�t>�9�C�*�c<Y���4mso,c=�&�@:����= M�꼴ׯH{�,ON�M4UJ�&�4؀4�`�M�7����k-Me��H�/�U����W��ų쾾��-˫-9�`�Bk�v:s����V ��"�.�P��/^���ܑ�Q�6�m͑	%�E�Ҷ��ee�ٗ�q�k�UxR�ґ���8�M� 2?��z�	o<�2P��C�[UWN�vw['��Zm���Ը��_��u�`:m�=���s���+W�,w?��ʊ\8���瀄�o�ʯ�b��7�b�n(���Z�1W���[Z9��q���pG*M��Y\�ﯝ���a=<B��&�3*�ͳ���;"*ؐ��=��@���޾{���-1^��6dm��"��΃��17�Lʄ!J˿�^2�A�py#x�u�1O'�␭���bI�C��h��>�r.Z��78�!6�Z��J|ż'S����ʗ�3g^�z�3�@�x��8ͱgN��	��d	��T���^]Rγ��/ss��p`�;.@!�ǔK�/#���+������w�����
���;oH[��յ@VE늮�&��s��Ӂ��X�t��&aUP'�ci5kf��bN�vk~{I�N|Ã@����`u����8`,�Z�M\lk��b2-<y���x��):���ǭ ����������!  ����q[�	���Ǵ���0A�C�+-X�����徖�3�C�e��:P�X[�g����g)��z�#�=���`�p���@*�jUjF(�x!��W(G�bGZ��N�22�:]_{�����I�^�Y��a��v���z0���r*I���<��<>>��E^�6�Nɥ�fE�����_L���ז"����x����s�\�;�M�#)q���� J��{�+���N˞Tip��!��Jܕ�u̥m	A����WS���#�k����sj5�kb��bA���L1#;�$Y��(x��(^=ӟ'�B��{��7��|U�<��\�G
vt�Wur^L��t�)hȻ-�to�*��w��`wgS�6�U:H1z����g����#���\�.]d՝�CjU!j�VrFՋx�!T�ˆ�SVۧܜ�����e鞌~����.���h%�F�P��Ӳ��"�&�T�#y���e^�>Ӑz�^ۧ�{A^y��SԘf_���M��{�Y�?���N� �x$[{cV���kȞ��1 m%cy�`�R������Y6����I�H;��,;�~-�U������C7�L�p3�f� <p0=�9NT�,�����¹zI:�r���{w��˵��3��bՆ�+ ���,5�P��/s�Iq9� &�!4<ONN� z��Ah�:�4w���S)�2N��A�w�J���3ZeŔ����2A%C� �3�^��T�TpXo��7�J��t]0���U� I����0��	@�x��'�[��6'B��k:w�	vNM���5�K�CO�I��j�Zw�z����g��F/6�z$ �XVD<꺷p�Q���R�7���;��~�eo��υC��^c� �G�����B�H�`�q4S
�Y��x�+@�ڣ�5�bB��H���J�o>Y}D�<�iF��4�F3����X�!t8-���?�����T:��d)g��q�\`,-#*R��,BhJѺ߾����Ŗr=�l�yZ2%�C]�]�c*��z_؟��}F7ԎT[& �f){�)�B? #���g�ҩ��k;�v��i4)���N�X�W���h�u$f�t�@�F�)���}�ܫ�
��q�4�����c�ٞ�P��p�H�y�ā��%O�� �p�"@�Y�7��ʰn�_�N����y������h|̆�����|�4��`��lK�f�
�b���IC�3�6�'�tM�<�)ƈC����!R4�X�E�*P�iԅ����ˁÈR����c��u������Weg��l���)�36�X���3���`�6���?�����^"=�g����*���r��Uy����O��C�R�2���5'��x�=���{i���-)5wr�⪥������6����H~��*��J�=�<��S����i���{�L���F%��}�=YY��3:�`��	�"�U�M���}h�~��pF��_��dA=���W \�.��5E�����ؐ�0z��L���H�!s��2�^��7x�c
0�����5�$�%���^D��i3�hx�xkG6���駟�'�\H_dya�F��>���~S^{�M��;K̭;K���eh!�r�����)�9�V�CϽ���+�R|+�SF��B\��F	Á�������Ο%��b��?���&pB��J^����*�����Na��>KkUø�&"F���~ז���y Į�)a��>��@j� ��Y�<OnU	� �`��-��N��N��a�Q�T�a��l ��
<.ra*������U�wYg(�d���c����F[@�&9�Z	�l<:��B�����?�_�벴ey���yz"�ޜ���'aQ�:�(x/�_�؃�j���m�g��w��0_�4t=f�n�  ������,߬ �TkR�j��~vC����X��kTٰ���u�$U��{i�n�hu0��*������גΫ��c�P�|4�6%D:;�Ԁq0#eM�A_���t�p!��c�5�$�;w������˧�?b��Vp��$��i��؟>mB��3�\���i��P�V���i#�����-XE4����}mQ�-Q��S����/��Gn�~+�_�h���*u#�fa�e�4*\�爞�r*��)�X7s. �g�-�T	��u�����~�9�1⒤P��9���r-"/�����ӱ�1Ҫ!�[i�Ʌ�OK�hOj�E���dS��_�8+_����\��{��Y��?���c�n��#�����o�/�ܸ-��j�����_��3�t�T� ���Vg��@� ��LB滨̓�j\r�~��*,�Γ�NBRH��q5̌�c���+�����C[i��S����;�X�5j||�ۿ,�,��',�~vü���lo=��yZ.�?+}pM�}�%�k����o$�?����'��J������(4�B:��zxP4�J��	��Ƈi��|��aȂFl��4�@a�t������������ˊjW��f"�Hݒ�
Lnݹ-����5^�N�V0��~��]6�c��Y�A�R}��g.'iY�sA���\�Nl<y��a=qŨ��b'�I��������i����T���d����m�8��|(	%�f#�����{�������`c"ꁯ��o˽h������T��NL�ظ땂TIn�ǔ���Lu����ʠRF��8�z�p
��1*>`��D%����g�R�OCO��W�)<'����;�+�=d�
�25��X�><�uT�>��W_��,'/?�|M���]�(���ʸ�)�>^�?�2��}8l��> +�,�C[��	<%���S��F��ë�:'I� 7F)#����ԇ�i�����;�`����r�_GRG#<�ն�W��d��Pmϩ�i��T��ľ�Gl=ޖqeh�I[�Ӗ��Ѷ"�����p s�8���)�ZJ���&%YR�?��[o������� �=
R!�C�
���a�we?��lE#;��VS�"�q���ċ�d���A.�8�Dd6R����K�7�mA�]��<���D��U���^������|_(xM٤���E�ЎJ 7O�k��Ф����z�2'�k��p������D�qj��Ի8#�t��5���a�r������>8��NC�O_�g�}�~�l>|S~�/������*o��<��l�q��LM!22Nɧ���@�x(uW�ɋy�����_Q�\�����lW��r�3g�l��*�@��%�0��9`\'�V��%*ON�W�QI��z�q]<xy�΂��pE��#��>7$�ր�[�NhM����tIU냃#���=��VJ�����?BoKk������7��-��?�?u��əs(�D�r���S��H��&�R¶�F�J��X�U%&�Í6-��*	E�Ղ�,iE
C\��/�&����.{�\8�y]�-�v�ݺsO�wwX�d�@[�)�l�����õh�6h<�$0�22��4j%?@��R��Τ�N��bފ��	{n0��x���V�'��=j=��X��
�� m��՜g�x���V�Z��t2)���s⌍���n�4z��0���Q
?�˯��ߒ���쫧�l��;< X�9��GzJ�����4D����R��iM���An��0v�a�� 9�oZe�a�����`����Z���#Ӌ���c�>h�H(ϳ��� ����O�v������wA�8,�}��yw>~�E6P{���4ut����v�7 @�Z6�?GU�F�bN�{�m!�z��B�M0�`�VA��a�v�w�g25�/�g�v�u��e��)@�1d���Y\ې�F���82ٴ��7�8��s�H���M��k�xL#DY���cS�Ł`��r�3��5��Z�z�;*z��Ha�|�KY��i������\��������_'�]��Ǳ�U��+x6 1�Pp;ܪ[7o'k�Յh�ژ�gm�Ԣ�G0�l��Z-��Z�a,�s� \p܂M���a ���jZ�}T� |4ԝX%|+8HZ���rs��A�G�gt8��e�Ͷ�:�������My��O$���������0������_�� �j�C:��/U�1��p:Nd��iYY� I]��=]WCut�� (�աk�N�얮Z
�v;)E]9�Q>�_�T��\_(P��ZVI�E�z� j�Pb�2��Sg���+rot ����;:��C��z$;�)�����[Z�����dme�]�y����)y����у����җ�ҷum���[.�4��6b� �IA2�S;�P@ϥ�pQ�S�D�,[c�!&��c��b$/���𦿃��7)�M�d��p���tѬ��ʺ��C�%A��.H9�0���2=R�&��qc)')�9��8�]��F�SEn0\�)>�<��q���gǠ��=M-��(��j��L��u�m*$P�H^��O�|���,�t�{{�2<S)��l�1�q:T�!r1�,�|��Y&ݞ�k����DM����H�\|L�uh4�h!�MM]�P�D��/�����h��r�X6��xV�a���X��4u�/)�'�?���$-�+*�!7��:zL�ܪ��P�5�ܗ���������Rԟ�;�����z��s�ML��h]�!���0��j�{@�>p�4��S��`HQ���ق��Rf���Y55k�W�����ԇ=Y�d�����vv��,)�������q�Q�~�I�~yy�k�;�[���~���M�Ա`i$8�&:�K:?
�9
ɛHWgC��K=���a��!eVI��sY�f`�@���d?1E�N>[.�p|�Ǽ*_���x�ǅ���ѿGY���֋��~?\; ����#_f����&N�i����}Ӝ!؄�D���0%&��B%� _��BjA�X%C��,�gN[�W�B!p@��ҍ�@���&�t��s�� 󠷯 e*�J./~����s�?�C��￮�z,�}�@�����#�'R�����57;r�'��3/KEA�����\U���so�
�-S�
ׁ6�N����s��~�xQSE4�I�~T�3��/��5P-p&x㎸r�.TB�^=7�ڭ��pI���'��m�S�CE����m,�v�dp"�X�>���5n�a��΢�w�#O�e�y(����r��3�s#:Tc�v�UEBG��ZMHUg��l�ˬ�Eix��FF�Hq�~�Ģ�q�Y�Z�Ί#�q�͇��u<��ȲbE��t:���z�$�[z���oo�0Lh ���O�r����� 
��ٗ!!�?��z�V����ʣ��D��t6��Q���pO�9%�L=!x�V���D^�����������U�PM�����	B���ɱF ���|L�DY6<�����ME(<x�hⅰ�����/�2�)�����\٠^JP~�C	�o���F��E9��x}m���Myxqy��������7��}�{V��� 24RھU����CHs/�|�l�?t���O�c'l�a@L�Z�D�s��/p@R ��c���R�1<��:H,��Z(N܎H�5V��&%�
s��y����2j�l v�E�Y�`ցQ�����I�}�{��"�u� �'Vz
�9t^�q��~=N\wz�u�>�u�Y]���0���f�<scDiDVh?���S=�O���+�
��(��W�VS4�T0�G����h�k�V��+�5�Ft�:���/���>o� ��F�ϋ,i���kN:.�:��n/Njc��Ui�-8R�\M}ޫ3 �Ӌi�&�_U��,!��=o\�iYH��E��@$��Z�g����	�B2���@0�a8�in�8UK�Xyxh��TeE��"���$��^oG�����xZ^��/ɣ��ʍ�ߓJkU;z��q�����?�.ͥ]Y?{�|��ܲ:PM��84{��#V��3�]��!mE읕��$�M�[��������B�J�;NG��1��t�J�q�F�Rʐt"�R!z馇���$|��u�+��Q��G��a�7*#�{�N�a�,�7U�ݗ~�<|$���+j�W$9T��Y^���0�V7͓1Ks퐎�s+�g�5ka���=vĒO���#Ah|�_7���d��E(^��>��c��"� �]m���j��м.~t]MjM��z��R����4<u56��`��
ý,[� ������Ɯ�> �SC��s�p�[(<犂%�D��h��041>�4�i�)#�̲����~�;��uW�bhdTS���j����4xč�9�/�(�F4V��V���5B�D�P^��A��v��0��Gh��K�L[��X�b{q���33���օG"�J����.o)@�'����ݱ��t]�7 �
� �zATx�����	�+��y��ey��E���,D4Ľ����1;��ӆ�Չ�
����^?�����c���ְO��ӈ@�p<>��YO�<p���8?�(Tuq�����`�s�{@�j��:ӹ�X�2�M:4WF9��1��y�B�[_�A
&��2�4Ta���*91�55a@TV��@��1� /�߈�`~�B����PLO��sM[��/"�]�Pƃ�6+�H�u�=�LSY�,J:ߒ��,:w/^��߅����\a��~T_?ct�Ru=ܿ{��|ii��3��R�Bm��҇�z�Q��^�k�W_}Y6�W��;��-�ӹǳ���(�8P��@�w��� @�|S�~��~O���F�B��d�R$�Z=T݅6�ECT��O���^H9{��"�_6�5pp��x��)� л
}����~�I�L��!�V#"a�ci�.J��x��i:$PI�2�;,i U�0�����2t	\<R������A�(o�ñؑ��k���8��z2%��O�ƩBt{�����[N	�� ���9��u�S�~~�����8�vF�|O�?�Ǐ�Ʉ�F���	���Yi�/���l\z���ݣc}���耆h�;vF�0���ِ1���|Wm�3�V�A냕��!��O\_(P��զ�I6։�yHB���{�LN7D�a������I�uK.�4�A��},��=]�-���{�&ɲ�:��{�f�^�Yk���{�&6b#�)Iq�Hm��4ccF����@��F M��(��PI� 	��@���ꪮ��rό=�-s����݈�&�m�KdufF�[�u?�~�xӿG�G54�D�6g�wFǲ�ݕ[�B�8�y���jzn��Ʋw�ev"��dT9�x��"[u�qٗ���VAE�ف�8��
�3��L�Z!+^��RcO����NG�H����0R�ѩj�@�i~�ɯ�#��_��T�l4}��,}���n�(�ث���ӹ��f��V���:��� T��z}��J�VY2�#��>��F��|ԅsg�ᑇPk�i��g�J��B���R�*�8����*��J9�آp%��%`2�x��F��"ё�n|8I���N�v���רI���n��h�s��w8���o]�r���[�w�ܡV���=�@�:�1,�L�5��'4<�A���nz�=��0)k� �6��������bWш�f�o�1�1چ��j
DLa�46�u[��[;�H5����EY� ��-�7�B(�G�o3�Y�ٚ�y�g��ά���I�I��, �/���P�K�Q���j�DxhvM#��G��P_p�E��2ހ� '1�:�{cͪ��I"�|�ޯ��go����S�:44)לeXZ����}����E�c�1^#�{�\5t9Ps�=�2���V�M� ��ݯ������>'_����lc�VI	�|�y���l��1�Þ��Y{��{�e{o���#ڤH��Z�J���YÁ��������4�ǁ�V�5ʂD��v*�DUGK�+���a:�^<���J -�������R5g�,?C�+�6 8L\���O�ɘR�#T�%���v93t�7QB~�dq�Rk�y�qy���A�T�� 0���������zA�k��E\Oꫪ��J��'��kͩ�,��`��	���E�P��*hp���	�o=��R�/�p56IF��ǅ��'��~��l߿#w߿*�woHz�6e'�%%���)!q0v7?ZXs�uY�/<.���l�����*�(�Ha=V��LA�.
��(�f�Go�pS��J��_�����'�)R��Z��<��˚~;ZbE�MB��D��Π)�)g��4T2�h#�a�Y��9!J����jY&���9�{K��=988b���k�qP��d�33:a_�Ӻ��)�n�P��ޫ�.*9���"뢪O���g��mݧ���������3,] M;s�:@��3�7>�����J�a%C���N���)^��A�q�VU�7�N\́B�Oہ�fR�5B���Y�h@>����X"����\T5(E�G'����³�S�;����3���������r���lc���`썎:\]?���Wi�P�#\a�`��~	�]�1����K�^����+�6K�Jnm��EV ��g?��|����������n]�9*�l�U{W[�c:���gAL�_AB/�-I����H�4h�!y��$�2&����"�D�ma]�V��1)j�9/`���l+[s���`�&�ο�^�d�(���h�9��v�k{Ǫ��t���ɫ���[S���KA<��wZ�g�Y��^��z̅;�+���L�̋��\���S�EfTl��U��Β&2�k�+C>Ϝ9���'���%�$�]ȩ5��s��S�l�;p�z&Q�3!�2�3�h�>�R��)�xQ�j��}��/��ϴ=^�������w��v��P�G�'�djc�Z���}:,���^^����_�*P��LG�3��S��bgjY�O���ޖKM�����v~6�c���vk���C3f�6c�Lr�J�tq�8�݂�'E�Dy�Ɍ	#g��S?>� �$x�B�,����ZX��Sgeo�9ν2�I>���O�,���{RN�:#Kk��3O Q�Pf��HP��fLN�w��x�%����E�5�H�`�bD̰G�c⣯\e���5��Sx��V�Z�Q������)ZO�Y�F�1��G5�8bO�⋉��4�亨hx1-��OLwb�b��������(�s3�-��o
:t�9��� Ҍ�E�f�,m���Dfb콌�W�Y�����;��Mݻs��F�Bg�L�i�ϙ�ԑ��Lc�j�)�/}l2sN�	�#,^x��ZV0�r��9�Q �xaD4�����1��p�����s�`����*����?}Z޽~���LI{�v�)�<�ȃ{7�u.�V�� ������LN�����~A~���`1���M��~����k��!��A�����9�u�I��oy
{&�=�H�xFr4�t:�����M�5Q�p� �8-(ݙ|:����A����忔g�}V����S���;`�vk�U�7U��>��Uў*����,��mjj0Ë��yhXstp2w���4}������3u�K�.�e��yj)ˌ��0��� ��O��$A��Y����;��Z��}���?%/���<��޷��!��_�җ�G=��7W��zU׌�������5V�����CYE���H5���%xO{lS\�d�V��\~�	��O}�{���+��c�1����|�������AX.�=fgz������gf�9<R3���r�g1Qt�@�y4i-�d8��T���
�_��p��҄4�f�s�����ɭ�ތ#�.�Z�W���;�
A��p�BR���k�@�[��a�ͺ�u�<���$M����A)���� D�C����}�I��S�q�+)����Qe?9ʴ������B:�I�7\����ď�N�=\�YΙ��$�������r|pIv����@��-fЊ�^t���"��FY"�1�!u]���6ҪHM�lt���X&�Z�|���ƘKy�u���e��b��"A3��҆><',�D;2�񠜩���P.�X�Ԕ�7�R~�{<��A��:dw��x݄�(�3��[��uY�pJ�(/���6h�#������pި쾰�7�́g�
����Ӳ0CeѷD���V�0O�G_R2"�In[$�g����,h�h2�a�E�Mo�xQ\��~���
k��0�Ľ�P�B���k����Y���?O8��2rp��K�[o��e��3�0������sg婧���98��}�kJ7Z�>��$J��̈s�̧:*��upj�k+rѽ��a_�hk���j�L�$�����X[���I(1j7N�EADG���Q>���	�uu
�#�)�2{�[��3���U��v�
ī���b�1�,],��f�l�"C�ӭz��Q���֘�B�O��r:��.J-��0�	�:W����G�.v�TuD�_��r�ȁ�	�:�3Rw���$�������Y\^a��T��%R�D��#^x�7�cv��->+�rݷ���uuj=�a�{��яɧ>�i�.I����ܣ�hׯ_�;���� sY�x6�㳒������LkT�s[|_�{��8.K	�:$Î)H���3r��&�0��~���>̞���(�ߟ�C{�̠�^�̨h7O9V�%7�^s�J�[]O�,��]%�jG��{�}B��R��S�{{U�q_�߽�Nn,��Y5?���G��0����m���tidͽ�H�Á>��*��:�Z�+�M)4��Wn�b�l/��F5{t�qV�L(�@G����E[폯M���M�M����)/�Q��OE�3a�*�%Z'�zx������� 2��y^66Ϩ��TI0��\|��N�㭸�<����6�4l��S���k��k����bP��A\�i�`{����N�0�Zmև�P�t �E����#�Z⥆k�4�:��Om����׻[����.�*Q�����+����=:��ES��g0�Tr^�Fn�L	�$�`�_p�h��sh�I�3
R�3Y(�| !}>�rjj�YUz��De�I�Du��W����ڽC"��
a��iVB6w���:B0���h���2�V�Z̾�K�b��`<8�#R��@��
u�O��t" 2�(:򨡀n�pc�-�E�Ȫ������+���:%�۳.�s ȯ��R��"52&j���^07��>��Z�k�r����<-�όРy�;�` U�+�眤� �+M[c�*�V��	9,e�iV�fF4Y2>��rnagI��\�S�HY�L�K�=ߥ@�f�_��cme�ى��/v�剪�ʲ>�@��v(�B(�i��y*� )���1�I�Adt@�`���сD~t ������)��`�4��|� �^SЂ�GSvMHv������D��HY�YY)�ߨ2�J�䂹�-�۷o� �b�<7pWYK A�輘.v�w�=*�"Ѭ�J�͕W2ڌ sY��Y~`�)�պ�`�Ɠc�x�Q��W�QfR*����{��º2����(f;i�\=�g[
�1�4���Y0R���V����/3&v��t����6�~O GG�'�k�6
��F$�@Xp?h� T�<���e�,����KZ5frg�#V�s�POJ݇��,� ���v�Ab�e�5�#Z���ΟWG��B���W��q1qQ>pFV5LE�@�Z]QhJ��-�4�� ��o��؅���,D�bB2޿q!w���cY�t�UPT$|�D�����Rw��X����p���j�c��ǳ��k��ꢞ F9,�T���z��Ȼ^ptI̫H�Te�Ω)����|W[�1)3�tD�p(��N��g�iN),��d�l�#$PZ�Ĳ+R����%z���(���3 �������|�/WԽNMXv
�° Y-���&K�Ȭ�SG�Bղp�l�PS���g�"_�6�BՂ��p2�B�R޻�����*'O��H�[郩\�x1Le}�y�iJ�<�0�� �~Q��v�gn츯�4r&�Ƃ.xӬt�4\������b5Z��9��A�B4ئDD\iS�uP�����eE	�͑��%��F�sȢ��]q3�)�����2�����Wz��A0t�+��j�(���l<pYP��ȁ��_�;�"�"�w�lQ@J]�{�Q؀v��-6e�
>'�nO˱Ƈ�!òe��6���J3j���B� 3����D$G��bv��5�w����8�Bg����rxF�Ú�y�����5 ���n�C����`.���4UP�Y��ޅ��@F8*c�|+Q���>K(XQV�Vkr�"���X�%����b��.��j��B�桡���Z{�Eft�L'h� �lD��i;'����8X��%�C�:9S5�,��Xy�C~~���r�s�Ҩ)l�i�6�����%����Zq_Π��󠄼Cܻ��
X2��4��AkƩ�����g�"Ov՞�����Α� ��2RG���O�>�;�,>A)̴�n^(*3ˎxg�f�{A���~��	c�f�c]@m,yx�8�|	(�lE$L���A���mb+�j�{��\>N3���HkM�(
L��!Y�N��m�("r�%J��Ǖa�S�*]�Z���0+��b���	� �s��d�n�s��m�_����΂�$JH�K�Plo{�qC.z�2?�"�J1 (���� �Z�5����w�1�sA��_]]f����%H��pZ�.��%���0�$�{W�J�&~���F����L&ݜ.A�7���a�pp��@A������YgTC������N����Y���?dR ���O~R����Wkҁ�w�zYB�1��C��f������eF%��NY=��\s
��֎�05�\�qŕ
u*F#����_���R#��3F�(�-�鼐����� ���5�"c��L�p�[3�~�)����=3ot�Y�({Ɩ������uQXԫqƂ�~ �������A���T%��z��=�Dh���+d����f��ܸ�6"�Li7=Piʚ�C�O����Cՠ��ÑL����Zp;�bn@���C��0��)ޱW\�Iuu��C�>�W_�g��¡�h!���֒&s�2mͲ�$ed����s���e�Ds���O��@*��@�(����{��j�=�M�5c啰d����0g�$6�Ҵ�J�S�������5�U���_-�������b�rj�i�!`%V*�y�3p`���kv��?7���-��N�6.dpo,�+�
ZNܖ� ��$�	�}A �}�	��!��}���\I�{ VT��%��c ��	�L=� -��NW"m{��qѡ�,{�*�	0��d��˧?�q9w��4��oˤ��ܹ>�c�*P�Q�5Gq��di��6��N̪��
lݕ�_�EfNPsC�ͅ�t{��B� ��Z�|�nO8M׈wX�0�X\�d��}�q�"j�Έ��nM`�Aʹ(��ȃHG��.��:2��6���@uC���S[�E(2�K�x,躞:��2X۹��[^�~�hW�T�Lc�w\�E�3Ť�zlHN����2IŚ�4��3>=h�mU���h��(��F-�RϿ�˿,����_�F�-����s��<�ú7��p�y��ʌ�!+-����f(�f\��hz- �A��&ŚAd�nZez�YA4T�)S�> (@`mwg_�7���sU|y���w�,<�� $�Ug�	�D��J��s�����Uܹ�����-y4ɿ��ƉU�~��0�ܫ�[��_�{é']g��Z°=F�uy�7��x�Fݓ���ynR����$�˴�p�\U��h���FZ�Ro����H�U�P<ˬ������9KSڪ�m�3�z4�F.YT	��`_�V�l��Q \u��>XfДlm������R�fޱJ�A�x�:�)�A���ݞ:�|����U�Q����07��4�-!q2p�y(�#��/�rg��,@V��/x� �"�lh6��8XnU4��߽�>�G�i�(���u�ܽ����"}��Q� !�A4��zdQ1=�;�N�����L�Ym��dLp�`����9�ʄ`%��X����J P�M�7��(�r h8� ��5����cS'	a��aOc��	d�?����	�m�܍Sg�o� )�� �٬F�g�U�E�E��
�g�a�f�Z�[�N�J�
Ҭ����.��>A�'��Z�5c� �A�P�"�"��@�mTm��3�)��&gُs�Е���WM�"ΌHʊ�8�i������Μ'O��u&����	�Q��f�[��Μu�ۆ��<���8�����Tm�?���%���[\	��hvw=�ۑQ�"7�L�=F�(��p�T��9����źS_(�fO��E?���])KB���I����f� �z:�ͽ��c*I�|Z�$��j:�ژ嵕?�1���H������h7O�qɗ��cDƝ��S/nVh����{�8VuJf��ؓ��#�����l��t�θ��x; ��@�"O?�e�ѥ�
�����*�I�[�Ox���0��4:��JߗQ��^�+�Y�;;���P���F�>�28��ӭ�t�K��X^Y�UD�Ю^{��`����ɏ���ɚ�	��謏�俚��Q�Qj�ܽ}[R��fj����iQѨ� #��^���{����3O]aϟ��?��;��|ā�B�j;q_�a�lGF��t(7o�t`^��ڙ���CXnL2jD�Zf)�I��-���E�O��=��E�fhC.A�A��v�䘉�o���}+��gں�Ny��q��q���M��\,|�� x��Tm�Ձg�-��rt�ְ�����3���P�\��A�����"5NI}(���La��yw�j$�W�sZ�)�CCbr��:mi8��3%���U���?��S?Y��{���ڞ��˒�CvO�ޛ`���Hf;�w!h�P4p�i5�Ԟg�EG��j�(7��(ښU ����K�P.m�T�?fAb�yQ\fk�:5h��5F#��.ȍ��6P;�rP��A�l�ڑ�[�=�W��s�`Pg?r!P:}�����NL��N�_QaB�Ȇf�)�9���IX�� ��� �}�4�o�I���&o1�Xb�Y�$n��Q_:�eͰ����J<�]����@e���p0(&�ak<=lT?��P��$�E���\�$v FU;.�:���l�D:/q?Cd�GUDHH�A��5u����%ڼ"*�:\�)P�+ƅ��|���e�ma#�IO�Wn E�B)χ�Q��(J�ST���)L��iMp>���񞙨�މ�~�ﵥ2���a�j�Q6�2ҭ�rӔ0�'ȾA}�����IjIT��8�����/��?��|��\�X�o���\�x��Ϳ���N=}��4�B�ݎʨT�D{�9-��E��)�[��j_�`TI�,*�/\�<�G?���s@�'�����L���������F����������[D�1cB�S/F����ӧ�ҥK�!.� $����+���H���B�I����O����ԉ5y饗��guN�;�ޑk7o�O�?/��/��
D�ۈ���X �N�Rs��M��Z��F�%w����@� �D�k�Hأer�AM������N2F`"%ת真99�U���y���(��o+�ŕ����j��0�o��I��,�@lɥ��bdgy-�5
��w�l��.��% ��O<缤t"�i��.��4.ɻJ���s2�q=*���䉂|�������ɰ;f	*g[ADjI�\�
Tԧz�n�0ҌS�JA�H"���}��'D܉e���Y�Ʊv�寐�U��Wp 5�?�8���C�����yZ�>ˋY )�ȭ�#ʓ�硕��\��\%"HN�e�S/�g��*��� �;m�.�5���o�����sԦiMI��Nw]0����O���Ue��<L�e��7��_2��j� x"Xe*�v��%f_G]��h�oUg�{�WQ6v|e� S{�M.U���`B��J�Xo�g�Z�A(��ZQ�k _#w�T,�ei!��{B�)�C��z�ç�[u�����}�Y��4+���C*I܎��"AF؀QM)�c�&�,6I��T��P�*!\�����H�p
���4)�r#Dxo:5pPܼ�� 2�X���<�q&%�$�mUIR=%1��B۪���{�\o����(����X�lQ�a�0��k��䉓$~���l�g�S�s�z��:h��J�Q�\$Pfx<P���.���d�/S�� ���IH����K�)�5v��=���~���Q�f�^��}`��{�!TEC�:{m)��J++�`�޿l��ը�22��˗/�� �B�u����������ׂ{3v�9�sv���7S�aD�Ux0�A��Y>��3̄`s��b�;oF~ �yN
D�.�[ �O|BV�V�w�w����Ww�}�<�4�փ]u
C�1#��Fc
�Y�2�dLN=v�a{o�ٽIvB�������Q��$�I; ���!�k�!�����CUY³�0㥷S�i���m���7Kv��@�?g�/�g{m�`M������@E�9�{b�΃g]��`�����۲�*��lp8j�E��	p*�3[�RKJ9� ���@{�3̥��Sܛ�6!��m/��
�x��(*��xh�Uз�{ 
MfB9�����[�1�ـ��S+����B{�sQ%�Z	*h��L(���O�}�a���l`�	�U�+�;���Dn_p�|֒y�Μ�4��� \&J,<�Q��s@�G�n-�<F�� �
'�GU�F8�>c��s���,ohy�9���]BR��e�"�Ԃ�q(a@I߇n�I�����Ƃ�]`�5�T| 6�؇	�� ���l٭�}*�X���mn,�`�ɡQ(ό����Fہ�U���ҁ9b���J`�Jb#�J�U�X�7�y[n߽E��e�V2��=�Nz���2m��ɥ�����)�)N�� a5Cy���	�z�s�9�t�tv�1eMm�ɣ�0�{��/�0�����C{n�ݡS���*:��^SL61}(���t�ez�jnփh���Ajڦ�t�� 	�z[v�x�}c���d���Q�(0>o��Ԥ�+�!�q㊘!�yEAj�0����/G��+vspX��W�,���^��0-
N��(Pv�{��lOH�3g �Q�с����|:].'�O�O�0^K����׬�d��B��'�R�V��V�W��U:|+�(��C`!X�����D�����C-�z�
JAªLA ��Q��ΐB�2xJ���:[ �M�|�)ԛ���"2Ϩ�!��@�2�;9�>pF�Oq*��bm�UC9��m�3��2�o�/�ͮ���<-��r�M?�^~�M+ɒ��'I+�5S���]X>�$�A&E�������g��mi�a��{h̀���3� ~��ku�<Wdi��k "�Zh9Ql��5�3����6�Y�jlSu���%˓ ��� �qz��8V�7rN!�*��R�^�,�H�N��tHx�X�T�u�e�^�ƚ�ǦE+dTÀ� ��#ó��׀�i�Zm �v+�mG�#�Q8�fKC*s���,S�(�&څ�NGD�RuQ2�d������s�\_^�tjv�L�ү$�/�;���0V�3�cٜ��:	J�j۪��\(���D\�L[����,�F�E3��E�!B�$ 8�g[�JR?�ۢo���C3�bugiY��mD�l�J�-�1�ea�\pMƩL#���&�Sv��9S1���P�:�!�������/��� �J;��zDL�q����!��-�BӀ��=W	sHg���%�X�'�����f'�����@`JT˄�"�l����*zY#��A��܃E��ʚ�0���4c_K4�#ů�cL��(�Nd�dRՒ�SbsWj5eGcњ��u�tF�o��LҒ4��qRzK9�C�;t��v^ B��Pu8aQ�PM����C��ڎ-�saV�94h�ph�[\�޷]��>_����Gh����mU�	ya��~�rC�]��f��u�)�>G���T�#�z)8)�Ѹ$l�x�|�:�����c�߆���V�{<��#���o�'��ϕ���T���"�آ���T���>��瞖.ȍ�7��(9*P�U�xS�[��NF�	R��tb�UU��PMvDZ�G� 無����+nM������_;����=�|~t�u��]f	9�#�)���}	;2r�-�g\����g�_5R0]ԇ�v�yݖ1g��K���q��0 @��+�����~Wn߾/;�24A��n�͕f�.U#"ֶ���Z�I9L3b)�����c�=�ʰ�eХ�<�(� �;����:_��H��$�/e�[� pȢ)�k"m[�R�(�MY6+��ṮA�'��&��p�)�%�Q\�-\��{�R~�r���8ల�q�Bt�����ˎ���E�ț�H��q��ځz]4�lg��M�hs�-����k\�X�1�_(��e�phI�w��G�|�b�{n\�YT�1M<�.���T��G�K�P�>�O}��C�Uc3d����OR0�m�how�#:�Q���dF.�ٽ/����<�����UmoI���Պ�\�� ��d��e9y�32�F��4�=j.�8^%Jga��m=�yt�-rV4&�j!����B�v��q6���>zQ=��pɴ�w�#%o���2`�]�WS:��V�H���GVvA=x$C�nk�Kd�n$�� .1������{ �	RMu
]]�pp�gw�*����p@b�kj� fz�B������R�t�AJ�fA��w�DA���KS����z������@�gqe�L�S��G�uƾ;��̜GQՃ��xV�@
��
���0�4��<x/��f�(F��P�ޣ
h�CY���ع�05�<���?�^G=adR,+�����Z���;-Sd���@�d�G�,Q�,ە�;��x-S���'�� ��Y����;r������@�(hW�k:���L����=+�������s���O~�9�����;3l��cw�1��5����}���R[	�LG�`B����ɿ�~_����(Z��� ��Λ-�#U)��JN3���JU���
������|{����3����G�È�l7/�;-�)�;}dĆ���/�����T%�\|Z�Ӏ�KŻ��O����_�sVґ�A�ݡ�J�����m����"^�|y<p@�7�#(M��@a��Bji9�,Q�ؘR�H��3����t/�S�+��\��^�vHD#&Bc��V�L�	���7oߤ�k�	�ŏ4X_?9����l�VR��	ai�l������~V�B�����f�qT��
Rp!W�{G�w���s@����S-$��vI�v�)�23����H�����7rl�O�t�|x����K�J�0�PY�HI�<�r��h����(ҙ��v�K�h/	}*�vJ�N�ήl˸G���p霼��ge��)��GO5PC����d�wIW���ݾ'k����]�uJ���aS��k��S��<J��2�7Sד�W����[����Y�IT�� ��R>���wwv�Hr��I�������i���(GbuG��V���C �7Nȷ@���ޑ,/��!}ui���rNvum��.n�ߦ�
��-RݖC�b�T���1�C� ���AAJn��vh��'b��GDo��lf#�_0��s2m�^2���:�T�˖SS;5��ۧ!#���ϫlN��+�b)y���8���LA�j���W��}�@.���%Iك8~���1��T?{�X�m�`�=tZ��\��{�P��Ŏ�	����a_I�Ȭ�C��4B����I��4��B3���4d|&�A�{m�ׇ�
$�W|i��ν-�B��ײ3ᚬ{��^��<\����>�����k_}�M�98��3g�$� �OMDdh%���]�,����tM�(�̰��L�=���5��m�Y=d/0��p���Ag�̥(*�<H��i�&K^�g��keI}��z���t�3�M%�iJ<�:*߯�Ț�qS���4�m�x\$�C:�@�o=�B�ʵj�0�Ƚfg���σ�d�N����Q�Ybsw�e���~߻�ŎJ���2t� ��=;�bɨ����.�r1��iE�Y��Z�N(]�:L�X�AVfcK�d,*^�k�|��;�#��W������Q�+�)��n�/"�=�D��╊�$h{Ժ�#�����O�{v8ܥY�_�pK�.l�����"m�޾��C��1��ì2v_J��E��"󂕅]ey^&��<�����6n��DJB�*�vN���������FqZ#(!�֯-�����z������Xe������X�*�~��d˻{�d �V$�-=��7�I=������{��lݖ�o~G^���r��������HؕN�I�0��ֵJ�<��뚳	6OȖ����Ay��sġ���. ��(�hF$��d?���̑��������������p� ��r��`���,�� VA��Z�8�DKAI!�"�)Ȼo�&���$����qR2�I�<{^���,�<#��?)���FXv�g�/✤+vy�V����0���	�
JjC�+WUW0��W�!�0S�;c@7&�*��'��F#T!�o�z����1e6o��H�[��v"���հ-LB�@��=Q�$�&:�)�P���\ˤnQ��$4l��=��g��7�E���EC�H@���k��/����[y*-f،����VVa��ma�!�O#%Uc���ڲ���5�i�W`ũ�� a���m�kv��y��C_��%O]�D��ӛd��׿�unf}n�p~�:�i�8�t�"v�a�4�9�--�K&ɖ���y�m�}��H�v�#Y^]������s犑�&Ƅh~y���L*�G���t]� C0��XQ����@����?j��0piN���|2?��^�(��I����FC62�{Ӽ�����H���>�9A<",f�
����R���߇�6+�Ay��Ua�t�8|s��$��Amp�c/Z�ޛ�|8�C��w�"�r#�:8���<��o;[����֑���|>I�e�w����R�`8e��s��t�J�^���+@��ThMs�wYG���L�J�#؛���+;���;Fƚ�t{2hjv���x;���,�4����D�g��I�9x���l�����)�^A%���]����Q�V�qw�g�a�'�r�l6?{���|�	86I�D�e��&\Pڌ�d���
[7g��[T�	6���y=�8'H�l�BK�<�z�ys
�r�Np��[�C"��)�_#����#�,ص��Z��n��n��'��g������C�g� ��ޕo�,����$�Ky�Jc|(��-���g��_�E��7�#�o�w��%+˅�FC��Z��e��'��ߒ���������9�.�v��]��ɵUv��n�?Q�7R�
��ԯ�H=�O
a��V������3*�(ʲVL �U��&��!��t�$���j��.4E�;-i���r���d�3P�ђ�yg>����"6����ܾ}C�=�,��(+n���AP�t8v�3d778K'�12Qս��aG���t�D���RhM�6#��d���yG�$"fF�`q���9"�.J	YۜVp#*v��g�E{��	9 8��^lP!D��J>�:ᤚM��v���?#.JA6VW��G�a�d�(	KNaˣiv��,ml �:?�=-겣,-w��2:��f;b�d�r�dp^$3�䶂)�D�{���D�'2�rq0y;�%	D�,�06�m��J�>�$ص�^U�m�kk��G>*G;;r���?��_�S.���g���`���o�)���V*�����Vj#s�®��:��>��an�
���[�.1��[��๊��M��=)�|��jO��El���|D�x ]��I�U�Ҫ�h*)���|&�ds��a漫Qe��av2�r!8�!{�~$ �҈DX���,�Ԍ�$0�����\!�~�G]%��G�tw��֊N0��;��Nw��I���K<�*�Ԉ?�لB�M	�(S�="o�WW���Ǉ�mD�.RV��<ܓ	F��.=�&�r�����!��+p�H��|��#Q��GRi�X'�i� 4�6,ה$��Fi'N���ٳ�,�פ�Ę֕�����%�k�4SU�����ʯ��ԫ6���g�(���$YV]�q�nPYދ���磑����#)T��(8.Y>�!;y��l�Kj�YAo�j ��wA������?��,�s�t~C�~���zK6V6���ݾ)��o}YVV7�o���lm0����1	ߓi����-��\��s"��+r8Hyz�)K�I�I��@��R��*�q����>�K?!dZ�HL�XT���������i2����~�����ٹwK�AӘ��ޑ�g���ɓr�r�}���[Ｍ�ݰ��]������i���3K.Z�6�T+�M���d��/��@��D�8�7*�y�.T�8�\lcmR޹�ک7�.8;㓐0)A�iF�J7Vug��F��9��?� ��d9�OyY�7 "��9J$���K��4s�/J��!�03g%�g�W��ܘ3b����´130q2󳢘��Ɖ�/�^v[r2�T @�C_���R���2���Ԍɫ��U�}�M��7O-�SO=�<���唣n_vv�hd�ݮ�OR��>��ǀ�Y�{��rkK�חeí�{������5��)x�D���!'V���
�(jBl��*��N�2�S��OK�#F���^�p��l�)~��aV�����ua@z�oCp��[��
��䖔�H����e��*�6c��2؝$�oS���2��ٽ�#[$�j)�q�������)ՉQjY�@@���y�y���oR�t8}O3a�L�c'�l7����؂2��o:[׌Hr>s�\r_���u�e��K(�f����I�vI����֡�q�!�ya V82��� ȗh�,�k�;����=O�|�>h1R�q���+��U"����Jx�z����K��=�������t& 5�1_���ףH�V��5���]� ۛI�Y��Z�Pu�b��5S6�9 ���_!�+�Vu�T�w�����[7���R��?'O=���+̎�w���������/~�������{��/�?L̜v�(Q��ߓ��{���'���[�l�3�d�^��*x�!%@�A�1�$���C*�DQOIs�,���O���;n����,���[W��W_�l�6�pK9urI.�?�L� ʊ,-`xl�T:�ι�� ����������ҮˉSg$�<���]��;�	J�插�*?��>Ͻِ�|s�������x���4"�YO4�0��C���iɖQ���T�:��MVN����8�����gk���ɲ�#b.�s��f�f���a8`LTm���ZcHh�/���'��P� ��[�ÒPX���q��:8��w��?�Gn&ӏM��{�Tz�<�y!�,a�&h���D���,�)�XU7���S�<���L{�M���.��:'���ų��yt����;�H�}�޽;�n�fk5b�3`�D:@�j����|�%��x�����`��`&���uMT�J����"�5{��R}�e�f�\w�S=�|ް�`"��
�aX���Ͽ�}�Fo��q�xW�D徵��x�0�Y � _hqm����e39����P^-���F�F��:����/����F��>����_��q��)��ۓt8Ri�B�d�90a��RF�j�_���يz߭<���M��Dy*����'�F�t��,���!H�_�����^s�5�C�>���`��)Jݕ�zuH��k3�$�3�^���[�5 ��W�3b��3�9�Q�b]㜞`�X�By��<!��l6�2���2�,�<���8���`�3h���B�\�/�;2ܙd#u�ymfO(�L�iC;q-�ݛ�e��%����n����Ҋ����w����6�u��u�ݳ����)"�+'VX2�?�g3	����I�ɭ���c�����mY?��\޷�����HgoY�7T��3�U#����:>d��(N�!՚�֮�h��LO�!��碒�}�v�y���I��%�ci������8-�М�Xa�~���!y��'�����kNxM�L���P������ ~L�~%i���&>��Ԗ��SK6J*�)L^��GT�8�j�L�2MY�D��^��>Vq��+uZj]�bt���#����"�I$�I5N������蜌�xCM�e������m9,�����eC�
(e�Db6C$|������=Tzp���ԡ;o�߽[4���.d�~%??���F7�ul�Pӹ�a]$�B�����n�Q*E�"�L d�z����#Ӭ�3�Ww��w|()2z� \<N._��ɺ�!��ɻ�o�}���g�U(i͜�EBi�!���z�]!#?tY4�k)�����Z�� �H��"r?5Z���̊ʉ�gLf�C�M��n��:��̙HDi-RQF�{�^ee� �Ϡr(�י� �����5/���yUZ$KuBn�=pҠ-�� �3�D���6hgԛ-F�P�E�������.H���Hw -��XHTe��Q&3ת��l����|��E�s��;�Y6��X5k�Ɇ9Wl���"r�ܺ���o��o���ߔ�h�4O@��bV�hl�g�ug$j<O�G�*��s��H��wCf�� ����k5�3�a�sVhkw��$��Bv�d�ͅr��iP�+/�1yO��(s͉/?_E�3����m(��lw(�һ�b�F�r����Z"�ᑳI*w\�ƚQG;r#�p@�3̼�ʕ��#�w�:�R�+K���V2�[�n����_����|�F{���)y���/�@���'@
d9���t����O�������pIw��<غ-W���#���{.q�K��p ��o��Ҥ��#����!��qk�&-<Lj�Һj�lQ��@�(A�����w����$?| �%��``��XN���N3��������8��Yh��Skθ6���9�ˠ�i���H�nQ�4Ʋ��܂v�#nH,4Ri!���j��*���$$��2�'��'��uG���+���V��	��#%t"���#iϓ��������(�#���^�s���7�EQ��E�2Ά�zT#������8T5fҶ
?p���TYVe>`�up�x�<�P+��|t�#�d1#fF�R��{���ae�g����h��=nݾI���"���_��_y��A�B�C�:���}J7#����I��9�A��ǈH'��4����@��8�<��l���G�RK��]񻏼�1��_��v""\�X�����o���1�ڱ4���p���#��/�#�;�����r�@�8��q'�@ll��_��&����h���q�:;C����5`�":�|�Mk�<Ε[�g�Pb�g��s�p�TZ�E�G��#u�?5-A4��8�F+�x�>}�S���gϺk�%���3�{�>��L˓����Y*lh�T���ă�N���.�Hթq��D�L�	�g!�Q�l����\��ߓ��T-���"*�eY�ݮW�@X��/��+�,+{���g!��gX��� ������ġ�K�3�Jbh&�;fa�;�MXo�y�lF���L�:>��br �fJ���m��zA�2"i�Unb�����>p���|��e����_~�e�����`+��,�La�u���ͯ�:��aU�pM�:�k�F��:a�k�����9̀Z@0�|ڂ�d�����K�s��$(�����ͧ�Q���;2>ؑ�u���\<{Z���mݓW�_c���}������+O� ~�kt��/�md��O�����_���5��`[�� ��eg�<�����e��Av4�_����z�|��W�K�'	��u䗥�N.��Z>8�NI@�ήq�gr��@��|O�����m�em�!�?{QN�XcKo�.����tz��/axa�!�%9s�CG}y0�r�xJP��O|V6ϟ�QԒ��\��
R�:�����b9��9OT�X��*�C�P�#s��/O�2峢fu�0R�t��v�y;~��-N�8��j��q�4Ԉ#�j��)��j���ŧ�� z�H3�1�[w����D���A� >����~��ރ� G5p����TQo������[	�"��5�������B/�-��gţ����; "M^ˡ��ᨯ�|�!����A 6���*�-)�͑x����`붦��C���0�	�A�0��;Y,c�3=�ʑ��֦������������7�s.�����.º��e^^��H��l�E�L2�^�R��Z�p �tB�sP���� _���bd_8����o����7�����-ק.������٬��R�c~}�gXv<�#g������N8C��i1(�t��o���*�~���|����{�x�d<k�[�D����pʈ�yr-�AOY_�FԮ���}��N�����Wk)�d���-4�ʽ�{�hH��t�Y��~z�[����q?o!�r_�%��?�������7�s?�_���/����|Gn:g�I�����sI�;O���{�|B>�Lm^��do����HJ�(;��,�د+?�_*2�wJ.���HΜ9G���>�9
$��3�������6� d�բm��LY�����L�����٭V���(4� Kޓ��"�`��$��ۻ����]����}�.���b��@]aĽ�n�}99f�	���FD��Ŏ\vk��mם��ݹO9��P��~n�:'��M쑨P˄*(%>��eYq�g8�{���޶ĺ���a`f�aY�j�*/EGx�xH�C���q|�@��hf�K��dN{*���E�T�`�Chhܓ���l�����e�ݐ�:7§~�Eg�Oru\��s��tn޺%�5��C����~���eՁ�f�9t}J~��?+�ؐ��g�|�/Wo}�=�%9�+��y@��I�6��F��S�1�~�1�����-иܜb.�(|J1gve hm �p�}��%�'�Ep�%�16@��I�L�mɣ*j)<�Ύ�!����(U�mȯc�"ĩPö:�MD����P�*�b����Ǩ7�2�!���R��,%�"#�C�?��q�o�R�}���ի-��!{���-�5��tJ(�BN��:*m	W�/=Y5�=k�+y��&�l�C�^�OJ.(���}��5w쾉�h�T[uw�v�>�~��j���7O��� ,wkۭGg��A��e4�2�v��m��1{�l�F��Yl�Ɖ�|������.����u���z�)�/�a��+��}̓7v����W<��Þ�<���9�	���C� ���� �G�k�8�ʗ��s>��q�/X!m_k�e�I�rj(aM�t�	�8~�#?OS��M���x����Ӊ���������8Y�(�F���Ҕ�M��3ͪ��3�^[泚X�LNn`�$2����%�i�M��+�?!�<�4�ǸWX�?��?�{��O�ݻw�7ޙᝄ�<<L��攅�pχ���0���9a:ۊ��2�u� ��?�_x��8���,�6��Ju�Q����ؓ�g�O���'�myR]wu��Rt�Ua��C���&"�`uyAj�ܽ%W�M�l�/Q]���{:�����)�l��L .p��V���
���v׳��$�>��<��9��w���iY^[�o�=µ#���Н�-�8�)�:Q��իr�ٙ�]t��ܸ�m~V�}�Dk�$e(1��	�DѶ��Ņ��ֹf9�Ë�R-��iO.�C[4kt|K�`=��l2������9�v([�ߗ|�w�3)��n^|\V��?��OP��杻Tx\[]w�¾!�nn��dʵ{8dk��Ӳ�ҧ?�1v�ˋ�FGΞ^������;r(��Y�߻���k�G���Q�':K�L�U��O���2U��\�d�(��t�q5���I�Fp�,u<`�����v��^������Z�S C"u��e̖`��Yp�H!�5:���Z9u�2)�/_�g[���,K��J����
��6����qLci5�Pi�\3E5|�E}_��D��֌H���
�ޭ�$Ӣj�5�+X�F��ެbn!U�[S쳂��w�a^F�y���%1���L߹��sv�DTAMY��x��DS�������w�bD���#��y��{G����΅f� n��Rm��[�
p���55t�#���{.��%��LE����3DUF�>Ð�lޱ��(_�T}���0�����h��ٔo�8��-���x�~�����vSpf����v��0�������7����3�<}VuB��#�d�i){��//�f>/D�,�\�Α
SD�L9>%U�;�Hɸv�x;���U(�zɝJ�����-���@�iy��cl��; upt�Rg�E�q������
�=�D�^
��L��:��Uv����s��ek�����d&q9q�J��Z��{eN��@O͗�‟���ml��7��B��c^,`ɼFV�*j��5�Gt���:Ǌ��DK�T�Ն�`D���Df.t�h��0V�I�Θew$�x��l�p�;F��,C4ҭ����r�剏,��<L�����|��g�B,�N�k�ꫯ2�x������8�*���7Bw��\�|@��
���Km;.p��7e����/��lɠ+��"����n>@���uX�w�c���*[3���Y���*P�[�"�����}k������I�8wCz����@j��=�svv�c.@4���7�:�<}�]:�ǅ��h���q�o�zK{#�x�Ef�\T��6��s���I���,���u�FMS�Ȫtn�l�o����L�ql���WNR0=�W����������[[������2�ĩ��1.Jgm�R�x8f��X[T!
c��՗~���B�Ѝ 3N[�3F�����R�R�-"2�:P�)Ө�^� &�5g��6�ؓ�p�G�v��3�]M����V�p�{���Eh�x�@�=�=D���.�NG�7�D��X	�iɬ�u4M��'��)�xT&�4�R2:ш+�*��6_��T󏥶Xy��Ԉ� c"�n}�����?���%Yr���/����s?���ډY�8%��������+SBČ��J���ٟ�Y�������s�
�cY�h�j�H����+�b�	�����΁WZM��$p�SmK&�0���'�av����x*���?��u��3�l��
�7<g�a�׳�zT��G�6����c�=��!� XO�f������=8�\���>9⾧]^ ����$:XT=����o>��#L,|�PMr�"|��+�ʅ���Et�a�"���1�=�����M�3V��r=h��̂�G��0S�AY�p]��=�j���02=�#���ܣ>#<��L����1�3y4k�x}�
��.8���K�kb����шر"h<t�-��<=x��1e��8e�]��[#u*�A�ϒJ����'���ζ\p���൲��`����W�����o崳� =����ko���*�����֎�'ڡ��|�+Ա�n#�o�����<8��6� -�^o��l&;伈�%�K@9ǻ�γ胒�x|�@��V�Y����[������t�e�����v�bcm�@a��������Qn8��n��Ϭ�p��������o�E$	��h�+3-� 0�c��T޹s(�n���*�]��:�GOk�w��x�-�}/�$ #�wya�[�m��ll�1g�W�-�9���;WֹQ@҃�?8��4Z���	� �^U�8t�Q%��ޡL��$n�Y�x� �e��������~���2K�R?����7~�7�ڵk�տ���N׹Θi�����C�"4fƏ�9��#��0Z�Y�25�]��ãJW�V3Z�h�T=�Ghלh7ȇ̺h54��3)��i�4)��@?����@q��;ը�;��U��<"�>Q�ɖf>`,�rk���SI��c�W(
�?�����9�|��tڑ	�(O�p@�9���O�K�ڴ�}�����$���(X���IF�Q%�_J�������B�9�>us��26���ZZ�R��֋�"fC,���j4�L�8�r�{�,3 d��=>:�^�Od
�y�Cfe�3:{攎�po�`2� �o���goo��ȧS%��ڰ���1&~�`$�4e�&_R��žݕjޑܸ}G���E@Y
Ο�@���.\B�z�<����}��S:����,��Ƀ�k<|�!H����Y����`M��i���9� �(#0*^�%� 
�Ą Ş �����Z�B {��Y���T�$-��a:���Ύ�9�}������:p��ި�q�7G����� ��xJ�؉�krtρ��b*��ǌ.��l_ۺ���cT�A�^DSO�(�67\�ږ��]�egG&�\���^ 7�������BK�|�WϞ9O0|����.��U�ZY~������f�>H�������W��m��-��|�:*���������f�3��%��d�E�K)�c	v�"���ª\�|^�~�9����D�T3f#@�Í@���u�ɻz�u��~&o�{U��[�ߐ�c���a���i�x������l?�O���Nj#m���c�9�zk	��noxUq�`Sz�~��3E/��v�t~ii�k���j#��`��P�X���Թ���8�['�W�hظQE���\B�n�6>��jLh�TYk�N_��9Z�i-h��/-����/83R�pkv�i�l`����Q��	���IS��0$ ���?�sY[^��%�sýh6�)`�tU��h��P7��*y+�2ǲ�nIf���1`[�����~��n�(���tw�.]�$+��r�!�ʹ��4���9���r8ȿ�7���St{��vJODڨ�0Z
�w�p��{��3X��p��q��KlfOi�����n�t6j���[��Q�a��W��t�G( �gYɭ�^��=��<Qª
�5��x�|�	��ţ����KxB�r��}���*[ֱ�ѱc�\�����E���9W��D۬�oAF�{����D���ߐ�V�-�H��zBm��1OGΦVHD�5��ߡ�IT�7��r��%�����r�#3/q���'����H+�k ,)�gX�����*幅"�cj
ť�:��2dH�5֖���PQ�1�K��_���U���f�}8�8�G$��-����'ݣ��̹�2<ܓ{���2�+�'E���3������N8�ŭgȷCt0�l�t<�~��r��%��c�; ���c9jk���6%:K�i�Μ��ׯ�!��O�%'m4qh��;2��qk��y.^a����n^K�d!���Haӊ��i3�G����C*�L#w�ڕ�#$C�$1쨁o�ȧ+�[�$�ȳ�7�~����KrrcMN�������_��9O=���Cna�����4<�.]P���9��!j�կSWVe����H^�vW�\���=�$�h¨<r`kW�wv��c+�� ����L���OUI7l	�(K?uv��6��a��{q1��}D����m�Ɛ�.&��9�B[#�e�����|*V`�-��B�6j����r��ӧ)��� � (p`l�0�,����2�0���%��< b����� [��qK2Z�X�}�e0�7O��{%��猭=�4����+���{�Y��:�t��J����m쇱a\�(t;<����+����[��������/}I.?��]4�� �����=EA�,A1I�	۲�� z�l�Π�t���풤��+�������ձ�$��|^e)��[6�;�G=��y��G��������~^�#�\51|�go�Kucυ�ף4Î�`_����Ih+ ���/ɽ�N<n�[�B9�Y�Z��_����pD�tPq�3�5o�+ ����$n����/-�/����nO�] 	�����㜺>��1�S|��ƃ1`B���e�Hf��K�Y�y&td��
9FH�`h$2�\�A?�������r�sBF�M�ࣀ^�%8�R�������7{���.�J���ݝ}���WOȅ�Vo�J��	�Ϝ=G��}� \"����m����w?Re��{��bM{�E���޺�5�j�r�<��G��ql�������]�Ʃ��l�����"1�A��l�<%��-/_fVv<Q�	Dy�S����7oܒ���8�&o��.g��t9{o01a�Zn;`�JY:t
�����|�6гˈ1��I��4k)?IӓyD2U���� -C�Z8w�WO���hY�#��҅�r��i��R�:��"�����5m?�Y��b:RN�SO^�"]���w\4�^>�E]L1�bV������}�Q�rH�E���N Zj����ʋ��j�vʇ�E�Q�S��b%�����h4�-�i�� ��Y�r,A�xT	�1�@$-'�덵1j��z��3=T�GU���vܔ^������|���gԉ�_|�_�i޼y[^����Q���G>]k�<)��J���~�Y�����a�`V�k�jx�ZD>�N�Z�+���yB��t�ɟ���������$��T"!�It�����Sz�",�� ��>���Y�y��J��?.��e=i������C-��ի����������%vF�א�G�sDJ4 ��E�"9Ӹ}[�3|�r"���L�~��ǲ�,t�^��44����8����Su�4�l�f~-��{�y����:�U�}���n�#\G� ��eKgʏ *�F��B�^3��'y��n%�}���𘳱�>j�C������˖��]�Ǆ�*��G�*�ǁ3֡� ������F'���%ᆳ�AC9w����p����l{��ɲ�Q�vM�Ĳ�e��G��6f%�3��>��;�]*�QQ�Xm����<�_?�y��5�3��6�1TU�"��׌�veV��Jϰ���29Z|a�D9H��� K�p�v�9V�,Ko���2)�/L����vN�Ȋl\�f��0��Փ���䄒t?�r!]�2K��w��m�A�\�����K�����~��p_wo�vӔ'�~����P���[��P���UM2�;���Vt�9$�l�"ǻ`�R�ǡ�	��b]�/A��#�9Y�4�-5Q�Ӗy�c���$��ۏ��������ƴ�!7:��F��1y�>���=��p�􊬭t��wޓ�n�����I�7�����������ӛ��@D�j/Í�޸��^&��-h]s?s�l�A���Bp
�?:t��vO�Ǻ�GM���Y%�>C˵�#)��\�I�ݣ��.��"� ��f	��޴I���w�9+k|��繛 $ EZ�DB4���a�#��Opx��`8�A2E�"%B@�@6	��ѯ<�y�js���Z���[�h�CG �b���̼y�9{\{-�s潌�����<�j�|jx�(�?�(AO{���hD0J���ٶ<��3���^�iv��2#�K����{�I�2ñ̏j��'�Gˎ��O��a|��g�&��,���]&|{� �ߑe^��o������'�w���쌼��+��s��^a�O2�r���D�L��M�D� ����E�VP,0	���Z�(�ch�F4��|�gЂV�w��]��?��3�):��
��~�&����Ϲ�Z�72=�!@�X dC@����H�0-�,凥�>���JT��}Q<¹=�5|K�G��oI���}P�I��#FP��:�j��`�ZT%�X�z��2:�T<�Js ��E�p�q��p�c�bS&dYh���&L����X���Y2��X[��P>�%7���q~��Rnw92��ġ�B)
� �T�� �5�~�Ĥ�`�ߣ��}�'��=���=U��o�T+�܀���qJ8�`�ȹ��u��X}�u�-���/�.G��	�g�A��J� �)q^��|%k���g!��My4�H��T�T��~굦�.#��Y<f �I!��0�z��qٹ�������/��Os<����������Y����y��������x��t�oh�ޒ��}��C��^Cզ�hIg~�6�AܐZ��8P''׀)�08X� O����>Od��ǧ���}�4([ES4�}H�
��[�̉�|b���=�A6u1����m��_��F|�{^̈Yd��Љ���G0���~Z�|�:؁�Fr���[�ਡ�����Y���H��(���2��$��d���W�\�U�G�?tX�Ŭt�v�Sb��3N�Ì�A�$5�AF��!�4�D��fE�77[�D=���U5ha�)3V�ܑ�!���`&�~Є�(BwM�~o�@rLL:��j��������n��`����e��䜠Ww����|��i�t�&�R~�Xw�D������v��p�鵛N�s�-��`F��g���op_����4������ǿ�qB+$�xaĩ3��_U6ܸ9�!ϭ��6�e�>���gI��X��
eJ��+q�0ǉ=����o��W��#�v]��Sg�5as!�@������`�ʹg���c�*2�,d�-u�����j��&����tձ�\L��d�7>e���_?��S�f��y���`�rAI��US:{-0�b ����K70��ܑ���Sq8�#�9c��3C��j��_g�m>�z��n7��;;�df �kɈWHgvo{�̦����L��������NX�OQ�@�M͔�I�I�aw[����+�ݭ�X�Dd�nO0�nE4xT5��?�������Vi9��)�2z�2��}uK?ƍ�9���?�zd%k��cL�4�
��*��ـ͉���m`�����u^�w�9I0�N>+������l�T���=�"��cVg'�4DIQ�0m�S5� %\��Tp�*-�'��d��a!����'����_�)7�ȿ��?�3���-���E���nL�,�4���>��� �>w{G��-5YU�R�m3�sGdn~������>��u�|�*a!�}Ž�:��Mz� �.X��{D	��x|���zE���p8�+�E����ǴE]7�8C�<�qZ�5�w�h���o��BGB��WV�������i�ҦS����GbmuGN�<��]�͒��Q������2�DHit�5��n
�~sΜ`��X,�Μ,;#��ϱ^ިj��)L	�/�M�;6r4)�gf@���5�9d|�A(J6���l�N׊�`Q�k���v����8��n�.J@A0	&�u�M��!�A��M�aPL�c���187 �!�v`<^�-;�8�`$D	�BD�����1��^����g�2Q\�G&��72sR�#��y��(��ŗ��a\����U��b<qdq8%���V��2B�lw��t����fX�q��,3�ݞ�`��0���(�s����J�-0�����I i��0�:X��m��&H6��r��'�����u���0���h���78��+�U�1`�t`�dLt���"� +u�ȘD�9^���y�����g��T�����o��<x�*���rou�%�j�I<K����v�?��r��W�B�+k�����M���������0����g�"4:��6f�D=�L�7oߒ?��/��^���Ӭ�6�5Ô|7w*�tt�F���LZ�M�N ���:$؛T���>:��^��C�D�}��C�/M��Jd�	��iq�@֪�c:hs$����YM��jT�b:���غ�j5��%���}��[�r�}��h�H���w�Y���>m��T�}5�˭#�-�X�]����ƠRp�UY=���Y�<� MX4���е�,�s�ff�ttVV�2hB�;�������=��1Hx������2_?$�NSz WD�Q/���e04�!����Ŗ�ʶ�����ן����D�J���o�}3��Ȍ\������r�#�3�йH�p^�V���jbZ�Ғ�峲��);�}�޻��7ޗ�����6�C�ߕ�yW?y��M��>X��&�di^�n��j��}�տ�X�o�ȡ�2��PhPؓJ��V��A��>�?3�},�Ǹ3�O@�awʪ��=����V>�@E3~��QH�2Ca��9+��*��#S�bǵ��m>��/ׯ��,�w�aڠә���Y�;L�����`�an^}b��رr��U���_ʝ���=5F�l���q��Q0�*w{#
�ud���N��;��u��	3�(�w0f[E�Y��HJ^��².��)�@|f�X�Ť��dD�Ը|���&����@U�}BPL�5|�xlKl�)kJ��>ր,t�H�^wnM)]`׈�6ۓz�xd���,�a"�@��$ �z`���(,�)������9�`��D�L���#�e�r��X �	%��b%L��P�@/�9����)G0A�����i��y^��!�1��������D&B�P�zB�u�y]���M`r�Z2p�;��#h��6�@ne��m��ZU6�ݕ?��'ǎ���m`���~�-	�P�u@~8UP`�����V`&�[�`S��1p���P�k4i�t�A�	%�5���v�veV��6�R�p��X���r�[n<�<���,>C��+O�x,�A�B����ϙV�5S�$�Z6��\���� ��l���I�5�`��֪�/]u*�l��{ο�ni"P����)�X���ޤao��4�}&�w�����Q���U�Q)$&� �{
̲XZ:��o��uM���RE!0Eun�������.����gc�@��2,���9wnޒ˗��r���)��s�&��� A&��'�1� �)�u;X%��}��?�W�<n���?\���"'<�����z�mVSQ]��G�������k����̒.r�"�=@1Z�8���Hpp�a�T\��#&Y@wpF�Ǟ|���V<�2��l��FJ�!�,����V-�P;�f;�_�5�t]�p�h��.C�2rW��X�c&�u�WGO<.]0�.�/{���4�ާ}]Ӌ�jT�;��Aez�m����^w�Вl�?zp�^�������!��)�#�T�g�Z���*��e;���X�'�o2� �~�vx��Q��>�"�h~S K��لIqZƽm����FsO�+����l�nw[����P� ژ��Cg�j-�����ڮ��l��������o^N�~��)�W�)���vC�F\2]� �2#B���jTF��Z�L��"eV@��w��`i�0�+2����Ž8�Fj�4Jw,�p�9�m�4iH�O��2����D����B�iH��AP��j8Vj^��@n:�� JȡNh�y��aZE���-�`�k�K`�1��"�R�(��s�V��aMi�ɤ����W;j(����?=�G>A��iy��/E�ՆV�:�h�F�b�����2L��`���
�b���U*C�I���I��1�쾺1ƾnZdպ1�v78Xd}Ǯ�	�&���qs�?p�j�2���O>mS[�A9<�N��_Ș�H��,��lƂ��X��_���}:D\;^2T�	�G�1������#����~4���؅�ӈ�l������s㧶B��b4�E�	�S��
�"�8S�HNqevV&�ɗ�r�90�4N�����*��9��{f���w :Z!�
X`��cD�a�k�����@�zU�B#8��
��BE����	pE8M�H�܂*�Y\ۖ-��l N8���SnkP������?���xȢ���	�*h�g��qpM�е:=M��T^W��i�  ��IDAT?\ƶ�:��9wj����.=�Vu���U��l�Sf��?Α��J�P#�*���ށ}� �X����
,M ��;�Q=�z�A�8;Ǡ���K��D��ڌ�bB�$l4�T�k���U}[�+��:��ܒh��#��t5���b�[X���Hw{U��+<#�L� q
P)��Րu=�UX�͖����#hZVkF��g�5#��<&s� !�(�CyC�I�>][wV��<����L�C���猦�'��jpeB�U\�֑��̽���Y��>���ƈ�;���5zC�wcm_�ߐV�.ˇ�u�q��r+tN�=#?�s�@.^�)o}�����`�4tA痤�����f��	d�a�@ u_���5J�T4n`�~��z˞���QNG��m���)�b�q��|i:���)J�����9���f%�8[�!	sc˔��Q6���H��^a�
%i�V=�cH�F�^�b�[]Y�N��έj����4Z�Ru�%� wHy��@!*c1|�l��YW���֩���q=�^G�IhY<5�
��e��X�hb�fa��s"5%�t�,��sDl(�� �S#m�{�2E&k����	���T�ƁU��Ĕ���k�$���IFM�Y����Cl�R���^T"c#�� ���$,+���CH>�dOW{0�Q�Jr�`��$�{?��r�M l�@���^�����Qg���:a>����ܹ������U�R˪�<6�	��t�|��{�$�+�A�Îi2f����4
�#�F��!�+E�O&Z��	�����z(����Ugh�̶-�0�er\FK @쿃�#�����!5���B��v//1�{��,Z��x��%����	���Bg����9�w��gԪ�mYK �L���"�YG��KH��NZ�FF���)w�l�㼁� N�Ջ	�1`��^�3���2<��G���+(��ma90y8.���޾�	0��r��e���@,�<�_�Ƈ����[��dc}}�Ԯ�R�vpR�A%�u��]��`�xp��vSF;#��AЧgV�>}ϮDYDHXA��;��q�Y@y�O���` �����D�#�4�����L���f���!�/��U��$Eø��
�T��9�c���v59Yݕ��]��N����1Y<zB*�YR�p]�4�/t�(�
G��������ɳN:?v5�gC>�G%
Su��CO\%ח��*�1�*F�@�O���l��fve�R��O�nFd���[���L��p��&L2�%^��o�;�L�Pi,�b7�3�(G��T�a��AƆbeuH�Y@� IqH�Ȁ��Z��U�ssGl_%�$&��[B�з+e$A��fhК�![Y_c���g��A8��6G�'�9k8�N�-'���x��
�v�,�q�m�z�}#� �f�z���:u��֮��_S.^�H <*ad"���XPa�Q8`Nt�� 4f�`*�+.���?sw�B�h�ː0PKo�����6QՍ<�R�&z8�d����u�ҕk�>��[���ש�q��}:��� [�D������D�/�䖑"08��T��c�aA����l.j�r������͵U�r�Iܪ͆45�FEqceW�>$O<���kFv��2��t��;G����ֆ��6��������'����'7�Z#�O�r/8�!���09}���}f�uF��&�qX9���+�<\A�e|�e��������wLe���Î�s�x�j��I�Z4�=�彾UXEvL�<�3�����ȍ_��W��j����g��Ǿt�Q �45�ρ{���������[o���!A"W�_w"5zL���Uh�����Qn����	P��z��%�:���<{��q��&+��6�X�85g��ro�	p��3�h���)��R�L�H����s�C��x���p[��G���<��S~�?�[�ԭ�c�@bL�1=����ؚ�UokE��1 N�4�X��sd��K�2�Y�X��g�Z��2P}����f��1⬠�Rk�JC;g��i�#�u��bR9j1}8B�Vǚ� iB�!a��|�:U$-}ϡ����g�cϿj�{�X�H��,Ā�>tMT�.�^�M����0�v�:+��>%���h�{TƅI���D��4� �Ί�f����|6�R�g.��ף����z���4���K=f�_&l��c=�`ћ[<*�kt4([43 n �±fC��=2)���] �x����)ݹ���h[F�F�==�qK�:*�O�� gD�P��`�7$�C��e؇,���1p���gr~C90b6ۤIh�~��m���п��	0����҄A�������>J��c�)�n%bF��v��b��۳�A{d̲!�s�=Gpӵw���~G���ox-�ssr����p��˄Q@��Z��Y�I�,5�L�{g!�ȁw	�¯`��H�U��K1DWg���6�. ��eKj����DWo�ۓ5͆�p=����k�1 }��&E-����Y���s��M -@�Tf���w�s��xZ��F����r��ay��W�٪���;r��5�ٔ��&G��xp�g���M��ю�����ϼ$��ܹs�׏ �Q���Jwo�(�Հ���M��N<�� �������u�'��9hp���9P�a�(0��ޠG�GRv�Y�N�MRL�����j:A�Ox-ʔ�e<ה���VT��q�(&\;8�h�X@4�#��SSg���*C���J�i�'�zEt��2��= ?���8�I���� ������D�i�{�V�ZӤ 2�8.�;[H����H'�߉�磀`ST�ڝ������Ͼ,���Pn^51���s{}wn<�٭	�*�jl@��m�	��@Y��0ܴ%y�<䐦�3_�~����� ����j>��ߓm�(�8 |������rЊq�����)87���Z&�Ǫ)ڄ�FS� �Sۋj
*xXo�����j�U��o���:$��2�>��U�g��F+}8�ODP�0�N� �x�Y��y�F�iO����@Z $�@dsw]��@Nj��|����w���kj��N
Q-��nw�[0��t極4��;-�����K��W%�F��Q��v/C�DF5���8�̦59���� _Q1P��B��3���ڍ̴�JC��=	k��xír��:)��E9�7����L�N"��À����TC����Q����*Ȱ���D�z4z�!$u��YY��CY���A!@�8q8r6k�>��4�s�(�1(�]6�H�e���`Vme}<
�Fv�I��Z)(�={Vf�fY&$�B78��P�/z�ʵI�n�3��,2��iꭈ������ޕ��9�w�X���o�̎��
?2z��C����/b���4�����%tR���9���Ϧ%[�!�u�ر��Ïl���@�┣�J�� �%����%D��MP��(.�*,O;��je"��S,�J��
�_���f!���i�:d�GW�)�� ��Kø7X�(;g ��X1=��{�Iͦ��Y9v�ܻ{]���r������ē'e��d�����z���?�����^�#�O�<}V��>.?��r��� ��t?'A���U[���q$=7td�L��
��R�Ǟe�`��8+t��69�A}�l��>��d�HK:Aa~���^ʪ�Y�r��w<�����WV�@�G98����]��Lފ�8��"k� p��C+�|�9K�j1`��#G���uc���3�����|�m��j�@�x�����9�}g�o ^P�������7��Q�"�OO�X�0�&-7c|�e~�#�쫿)�=��|�O�X�x��H���yԮb��s9�Ĥ�j{�|��������������ϔ���Z)���N�2?�쫋�@�al�wʯ�o�+*�T� �o�cM�e��J
	��͐S@��~�	:���eR5�	'� p��K��I#+]�T_o�`s`ڈQ���������5��e�J9��h�׉qs�01t�ĀF1v�*��{�/L�K���M[`�*Ξ�>����j�[r������'dgc]V�ݣ�ap'@�\U�>� ��4�]$�6�����ǹ;_p��MA�_S�*�|�A�N��i�X����ɏ��tǓI�8L�����@%���E���V���OΒ���J�v�%{�+2�/)4l$d��GB7��N�=E�Mz;}=d!i�%��>�('{NN�}F�!�;{$����ΰJ���d���B��{b���c~SR5���UF�ڱ��Y���� 078p�[���kT�93��m�15<�jV}w�&��l�# � ��&����]���޾����n?�Y� eQ�Eu�]��aO�P�kM#3�a�CD� c�9��I��q=������9���S�AN�¦���:���o@'~da�m)n��E�##�j��UgN���:B�����^�M�C�<��AU��8A�o�6�8���{h!��)  ��?�=C��V�A�C��S�Ԡ�����|�?��綼���Ïޗյ;��C9y�t����pm��~j�4��LE{���{�C���5y���r��iy����jh��@v6�%�Yr���{"���� "��8�1B�YE��,Ef#� �׈�B V���s
Rr ��U����<��q����A�w\�`&*)��@��fˣ��*&��/l�9훂1%H��2��e�r�.	]� ���X`��0 *7[`�&ax �(5�,H9r�t�|ݐ���u����w�μ��4A:&���|$���U�
V%��Rؔ�K�9��Z՜�n����U")����|�%'���E��m����1�B����I����6�>_�����Y=}��0�>i������~Xk#<T��by�d���5����>���rp��s�D��}M ㊝_�(�����\�Y,!��R	�p ~c�7Zt�׮_������-&�X���QL`��<X �D���"�
x҆gY"#�wq-}t��>��Q.��@L�0%F`�.�x.ưA��VUv�5�2[��_���ʂ�:K�t����c�/h�#�]\<�iF�v{��df~Q?w���ۻ{�@+�*�):}��gW¦T\���I�ȴG����-��^,���?>�@��V3٭�d�е,*����$=��1k��)�P���`KV�ߐ�Ֆ���ա�ە�����C�a��D��<h.�¡r��g�=���
���t��^�u|;c���%�6e�Z�w�I��N�ǀ�b8�a�����̀�eeW���á`#o3��C��=bG쳣���t�I<)m�ʅ����,��5��g�l=z�5��x�Ʃ��<��4p������a$`NR	���Sg<P�ȡ�F>@6Pm9��,��Tup���'��p#���f �vOӮv��j�N�+�ہD|�����`f�)����5���/�c/�gL�E����H��b�kS"@���[���j�.��G�8c�eA���ø�Q�>3��A����².9^2_S��*SW�E맩��W��Q��wߒ�|�5Y�\ՃH}�.�9��b���ki�?�^�z�}��vH��,u��z�@��\��+w���q9���4�r��\
r)�ċ����Se��K��h߸��2��-�j�J�oU��ޮ��~�s���O����}��w�YDª"dSQ�yP83pSTc8�+c���.�����{K�|�V*���+0>��؀�8���Hr�^�(��`�r��	�G�M�s�G��wߖ+W���� �[ǅ5:���p�#�q��l�n-��{�y9��$wnߔ����I`�x��Ѐ�9�C��S�[�#2��
x��{0������V�U'0�>�Ib�;(��%\T��%c��T�l��Q@�,��{ＥvuW*��{���	 #7��S�r���<;r�?��W������j�>�(1����V�Q��L=Q� <���!9u�Eno��|��Gr��u�$�tu�O��,3���d������R�+O<�~=)�.]��nߪ��-��5��B�l���� HN��;��"�l�e��@X?Xa"���¦V"�?�콰&�_��\	e8�z�������
��Z�/��pCGb�B@\kKG��F�1^�{/E��W�נݳ�zS�pD����Yt1��q`�F�!L
������Or�~o�>O]ϐ&�z�Q"��O���]Hu��+a�!�=�P�9{�����f^���Q�qmikDxh��f��d��k2��%u�>`�ƌn�Eiu��!�,,��V�Um�SNȸ�����4
	h����06�Kl�!�i4�E?�` �щ��a�p�S1�,+ݑ!4�C.������ab
�'P'̈���e%��S2�F�����w@$��B���R-a0�����8/dw@�4L,� �)��Z`�Q��(���#�3ebE4�o�#�����jD��* ���.H
7���������43��h�V�vw�@ FF�^1j}?���/���<��<ܕw��Юm���i<��q	l\�ʪ��k7yP�<�$_�Ν;V��4XJP�)�0�� �J��ɟG��&#c��!��
'�V�����:u�^��k�������Q��,Z�:�q�ƻ�Y��+ �����&�B�h��J�gd��ݭ�#S��ӏ���7�Ɏ~�$��S��"C;ʱz�!-���֍�z�	�9������Ω���~�K?+������9���g� >��C��P���I�)
���8�e��d��o�0s�F$<H�^~������S�c���E�L�әQGސťy�_��o�/��/�>�X���������1`ʈ���m��:�tں
8�q�G��>-3ton�XE�j�(ޣ ��!���H���![Q8�:]�(r��`:%)6����k�S�gH�$Ŕ�v4����}8k[�Hc��B�~��)��_��|ʑ#ˬ��|���_�����+����3�c/���hJA���)������]�0���+��a!4���SO=%/���<~���8y�{���^�ulh����c�Վ���7�2#؃t�t-����o��>��lYyR�ў�<0�����JlT����|���B�8a����NF��{X�>�S�vU�����	c�1t�	��x6Q2E�]�p�	n:��z��ߍ4io�R��)|m*�F���5�Ur�va U���F�_Q��#d�02r�l|��o��s�&?A���LQ�����#M+��~G��Ywq�ca���N5Sb7�Y�%ud�I���'do[z�-��#b`OQ��f{VaK7TM�F�c��.J�2��&�=	�
�:�9[dW���Q�8�v
��&g������X�=`	7c�8э7�$w�A��3��I��FVVu�Դ�A/<0�e���Eɸn�J��?�PL&��܏[�b"d(��FЩ��8d�,"������z�z�h��Qn"U��*E��E�$��j�^L݁����<���jH0*������в��縹�����1U#ۙ����_���x����w�/���-�� P�K_�Ey��geww����/�"�7-{z? ��k��k�5_�;��� �"2�b$;w�?��0�b�mq OjYi,+l�1'�^2Pg��l;4t�}��_VpZ��������m�_���A�f�����7��Ԭ����0� <���  ��t��ͤ���#������5s?!��eni��ܰo-L}���{�2ӎ}�����4�X���#�ij�9��8���3O�����"��@3@T��܊kIN9Z�O8��Ysyd����*)�$����2ۭ��`�Ң�\y�o�T֠��3g���7V5K^�V�&��Y�w!E}�l\�'S�0��:!��`U�7�u���V�`w�=�aw�xz��}�1��A*��(�~b��L�bU��p�a�}�X�<����W4Ъ��B�Pah�*��$���ٱ�Օ����|�-��쌼�*���8��}�{�޻�h��_��w������M�Ȅ����$^۫<��_i�[n� [����I�F�dQ%�Քٙ�O0t>pB���#� ^�P�cpvS^�q�I{�����1谭����+p�C��A!�F�uD��R���:�V��j�NLыT�#M��cr�AYzLe.)� U�]�jgb;A�}�꒗�v-G h��|\a0���Kw�Kft��0�S���G��]��i�a�뵶�;0�'27��ʛ�&���z��
�N�������S>�@�9�M�|��wF�G��0���f�F."=�M�;gg���HXO.Jt��ef�X#t�mc'� �g�fÂZ^�@v�[��X��\i2#�i��3���V@p���D݁�*I�R�3��� ��,E@ž��E���Ўq#��V"SF��Q�@���-̳��О��u�u2�*�M/��V���8ss�~$��e�JW�9��FK̈$�6�c���E��1��Ƚ���Rc|��z���le�Y	�x�g�yh�F��C���6&����S#�v��9z\?�P._��29����_�ӏ?!��뿑���T~~���瞗Uu��|����\�q�'H�j��c�-�h�٠��%&���^ᦩ���'ƣ��2'�}�������������}Gs^ZU��ߔj;�[8<+�vE΀{0*j`�֕����h��k?!Xkj Ziq-A���怙s�j�u��� 1[�}��M|P��X��HΤ��������,��H8�dTd�k� !�ue;��;�;����:Q}�GW<�(;.�O�L*'Ez ���xJ������_���Ԁ�V�N��8$���'�͐���a1	��w.XA�a���
�Ws��;�޹���K��;�{���yN1��L�mn���Sjd0��Z�g��J��y����d����e������7�)�/�ʪq 2�h-�C�?�I4e��Xn1=��a���,�T`x�-rcF��Mu-s�����WZ<��<	6!{�)�~��Sx/=��F��Z����!����z=_ ��yh5�d��f{p�ąw��U@�$Y���p�_x�ey��Y}]�P-�h`:�`c�3X�z;���R�L�J��
��V�zrv0p'v��$�`І*E��Z���Ɗl߻���^��A�%��/r���W��	epU͈���v-�f�&";�(��*��Mv�]�_\�������h�6�?����yak�^�ɟj�2\�,ٔ���rvo�&����	m9�w�����đ��&�񘀺�F��)H'�q<�I0j8LMk���d"���u�]�ݕ$���M"EVg%�TսZ���=�0(��[�vA���,�N�D�"�c� ��V�.ҮW�)�$PAkJi�� �՚��,>?�܉i����%\L����f:h�Xi�4��OA0䲙#�w�DZ�DS��V���%��}f+vh�� �̗�>>c�S#x��3�U���a&�l��������VJ`[<0�Y�m��U�銑���в���_�g�{A�ܺ���
3B�����z�]�y�~�������������ޗ��y�u	���ៜ���衣�%ua-���������C��ТҠ�ر#�ꫯ�/]�7�}GRLU�)Ij:�32��dh�i�7�W��h�k[�C2����"���^]_3���vF���.�JCj�V��A��~�0�(0~�l�25s2 ��`��a�!���9ރqw���J�d�ַ&A	���
s�M�͏����A�� &]���H*+8�ԙbX��[��>�1�z�J�p|��Μ�F�r�I3�#>A3�	HNUe�����!���Z�N��G�ݞf�3N3�ϒz�~���m�_ HA+6�Mwic#d$6"]{�e�y���kԐ�I� |@�����G����l7p\7b���������2�夗	"kǚ���J��T���hIz�lӔ�qyx���t�s2]{������;7�_T�Qak����5*��������2?Z��5��$vL�X�J%�n_~�ey�'����˔`�������4a{v�A(&� ��D\ \� �Qx�îU�2V2�[�U��l���β�C�i��6r��6�h�Ӄ���a�@���#�B�q��Sx�|0p /�6=Wl��vĻ���>1�m,�h�#�k_��X@��$�/J�I��p%+>����O5PA�+��h�kd[p�_&S*�3x��rだ����C��m̙�f�����@ �7��B"����K�`��������>#:�j��cDsLt�+(��ue�v�?q-��#p�$UM�Ц�Z�k�I�X-&��׊�!B����N�cnq�@[��w`��x��5�/`�e5�b�0;�+!�h���*U���	�mf��Ȍ��X`\�ԫ��0���N�5��
t�G��=0�ߓ:�(��,:LT���;�@���Vư����
���]fT�Ȳ�{a����̑� �ѯ��˗.K�� �I�,vk����>[q��^bZe��:Q�qJJd�f�
��/����|�_���m�t�;��h�f�sQo���j�0bN�n�{�;]`�`�gh�2#��+����ѩ@�Ծ�=���rh���.�ɞ�\Z���z��R�֠ _8`��{�1r	D��J�;�π�(@
�cJ�'w�ޓݝ}V"�`��l�	`��[KN��I�ҽ��
�p��LF�EPK���U:��SE&���g���Ԧ�V�Ij@�����P�#�xM��>zT�螬r���P `���B�����\K�_�51+.]��g�����\r#�HD�g�����[�B��g*q����&��B�Z����x�*�ް�9�%���8����o`����{��zq�Fz�ME��������O�
� p�Ol�)�!�Ē����I�������r��0�<uU~]�>��ARh��Z'��hg&%G�VƂ�HZ!�����o�V���1@mwf�W~J�IV�����_[���ߨܶ:h#������?�}?�38�}녬�BC/�8��/�v�s�ӄ��R�֏�k@�]�L[5�A
��A�DH��{���b�z/n�qTߪ��ƃ�q� �5�,0js��i�?T�oK��c=�ԆL��W�&	�C�6�Ir0*Ѻ,�v��{Y�	R�W�,&��lu�x����)�8�v<^;��aL�ئo�ɏ��8�������r����A�㜨ija ���c"� w����k9�W��]p3�����񎥢�[ᢎX=���Y��F���82l
FHI�T5�rS�/��W��A�z]��b�wRu�x��V9��4��172����o�YP��H:����+օ=y>g�Ц��_\:$3��̂�H���.W�\�az�XB�0��Hh�H�u��A6�U��ݓ��i�d�Z�Y(d���`�U2<T��E#�������
ȼ3 V�����<��sS�d�Y:1��k	��H�,Pq�V�ô*����58q�_[����6"�{
909�+�&��yN*0T�ɃQ�2���Z�e�ΖU��`�N�P��禫ƶG���L[z�=k!ۏ+�c������4G��Z�������;�/��h�6��A�|.Xs�������lt���Nc�?����T�=;�MI��!Z�I⸇ޘ�s�[���c���jAy ��K���i�������׆�}`$a�as��Bty0��g�)�T�
�u�L�����ڨsfx}b�0�����:�9ߞy	�wn�J�Opyl#�̄��t���AwT6��5b�����H��&����C��<TyܔɄO�Ah9)��]��o���zԞ)?�S?����ZUݱ�:�10��W>�����l㜭uh��s;���%��Uʹ�?$ �W�Q 9'lEhU�u}K��̑0�]�/����K���}����.x��C�׍[�L�ثh�By;��?6�TD��L���U	n�$��p�7�����y�G���Z��Zm����kB!�J���f\+/4,������[7��8���C��,�~BD	�Cßno��.����ev����!G+d�����b�U/"c��,��'���]���iAMT+3E�EvJPRww	xB�2v�z�Q2��ʛ�I0����
[Q�c$u�Y�[��֍]~��P۪��Y�A�d�[j,,���k1D�ˌW2�i@�vH#x8|�mVWWust� b�8���)�xf�1 ���N��F��α[N
�t�Y`�Wb>Ao�F���kR)9thQ~�|I^~�yI#f2��?��o���q�����d�=�|�Z�y�������ɾ��3�z#�j�M/`�b����2{_ffg��$����rkf�?ǿ��~�p0�Q������2���`{�I����\� �rzA�e�׾�-�8�-u>�#��--�k��6�
=fo5��ؑ#��������3,� \׀���;�j��+�vL���qB
���l�����'w����	]Bdmkk�er�ݺ~S>>���Y�޽���N�3_[۠X�4�rTI�U��Mk�5��c}� �dU%,&{7r�r�k-P$�J i1�9��	\˓uN�	+�0�f
��jV���?�ǯɹ>����� n��[�b#���*B�EE�������Zl"bdY��B�l���=��h�0��J	�l��0��HtI\A�z�imz/�q_0���)f�vf8�G�O\3B;�^u���QA<5�&{����v�**�;<X�H�}��g��p3ၽ[���}be6�Nq�ϓ�#�R��r�����}ES	�}pdmYC���\A��
[�����t�#�C�Ц"�W��-�V0�@���i@a�!�K*V��V{�����?8Ot��o+�*6ޓ�Zbl��*��ct�pL�Ǌ>g6�`pU�)_��p����D~"�MO���?~F�ҐX�#����s�'� �ah1����*e$4)[����^'�
���_�&�ײ��S�Z� M]T��a���끫���cE��D!E$��'�����(�n޺�n�B�gi�]�,4���`C��-N� �Bq���GX�@"��`HJj��"�T&�Z���ޗH3���::m�SEV��?�� �pY�vrW���<�~	#И-�"5c� �*bp�5k����"����H�����Z�������ˈ�ot���oP:`�oU��jtP�I��:�*ʅMи8Iz054���#�����דġA��*O ��	�aa�w��:�}5���_�/|�e��o~]><��#��|E^x��x鼼���rCbه:�c'N�o}���{�F2���@������p�Q����۴Q�c��/Qj|og��^d�/�t\N;.���WG:+�}�3���|�;ҙi��g��t�Y]��G�����ҩP�@i����^�ȠHR�*��}���ȝ9s��ëW.�8-��	�eg�#���b`QR��	������ c�@��[�0�`��#p�6l�qd���[��>w��ҨU�X	�i�s<\��c���+��N���l��n߸-�$��o'G�I��������Tۍ���T=�ήƑKR��L7	�F���������?TU� a��Ɂ�d2��\}���+#e�[%�m����l�N�5�'c%���hT"���]��Qu��;Q����D��(�#�v0��@�~��k�e����@!��0�9P6�WK�x�J�5z���� @�1Ҁ��yPf�����Q�Z)����"1K�=���uihp���>�.�jм����eM(��c�����ܸvA�^�"���P�Br9�C���o4)�YP���H�'L��T�S��`d����Ib?�56.XH�X���4���IS8-�"����0�aO��w���-����߾��X�Sj{0��ό�DLV�֦�9ɉ�A$N����!lx�y����AUuT�X=Fv9z�Xu�5�xPH�J�\��B"n�ИI�ъ#j������A,Y��}��H��̡S2�&�L���� �J��!��9}�~��I�bڇ�ت����� ��~֎KGmx<f�+$C���9��u����#d�O'�0ތ�����%�S|�Q	�q��o�4c��3�������W5k��ȹ�S7����C�~�`���y����+�g�	��gllh��!�GpA'�:m�������{p�ۥfơ�?�@��Ba!�eU7l��>`�:
�f�����l �f2�L�Ղ��iwZ<��L[��D��Щ����V��n(�1Wx��=��?��
c��Z�h7ڽvL���p�Ġ��ޫݗ�f���-�W#x��U��?�#��^����kRo5I(��e��Ufh����?�Q��|���<����:Q���E�&���H�����j0�<y���^���z���.��O�W��U��`�4װe����=�������q_�����[�9!V�)�����6�&�������W@�ڨ�̀юC��J��҂�I�U�z3�A���<��I]��Ƞ9P�/�zB��A
j�UQfF%A4�`�������j�X�q�H�<}y�Y�U�L�!�Q��>)����^�3�5�`����Ǆ�����3��롲���bR|�ҷ��b�V��!���L��IW�#~� �� �1�?�%aTj͆�%jU�g�@���=�u��ag�P:�6 �j���~j�5���m����\��� �BԈ�(��s7R똉����D��2��1Y�$�g	�#TqZ�h-TOl�kP�ْˬj���C�V+hw�ͧ�G���ĉ��M�j�o�j,��l!`�4�����׾��޹���ЎĨ+E2���xv�C�ETlpoPY#�����<�u�8�x�$L���ҙ�'�wgv����ഭή�X��!��q�ĵ�kU#��xm�₻�v�,	8e0�^"ۂ@��� ���}��E:S0��(�tMl�N�6Z_��� }@j���iN�bX @w���d����9͌&���j�/�xs�gZm�1����RЌ	���ή��pY�����s�WaI6vX������6Z��09��p�}�mV	k�CW�Il�"FM������]�v�՞%=�~�g{&:IlBӉ�A�1�[[~������o������ӨkC^�@v~�X�STz�aX�EM���Q�%��4g��ѓr��Y��ͅ,� �#f#��C*���2]lFlB,
��z�A��@�l�Sk����*��G�� ��z�th�
J�pd+�d�lf�¡�L�,H�"���� ��{G�)D���0�FF�I`{�y�!0�F���AA+g�j��V�f���m#0�F��3ص�F	-+���i!+7d�ʬȧ�v��,3�6*��&�j�u�]ɑ�*�����@�]�Ȓ;�Š�2zC�cP �ؐݽ}yV������>��ǯq��(y [P0p!�`��pR�ﰶ7n�p������~�������ϰ�����>���`�}�����6��4�P���؍u��MW�80�?iK��\�͘�K%Y;�����5���o�=��>zhٕ����j�O��qG�L
�v�@\����2B��w���H��_� 
T��YckW"�j��u���f#\�:#����
�;��丁�YR�3@@��T3*�,L6\����^o�YѠ3I���~�
����U�9��en�*$N�&��p�A�Ei��Yu	m��J��1x	�2K�>2����u�'�#�<׎�8���Ig�9%kyL[�t��r*vu��g5��x��е#��kA:,�&��ݍ�����L��:����ڄ�ri�����^�/u���� zB�hA�����}Y߹Ȫ��/���ԓŅ�:��T���Op���M%g��QR���i��Vǆ�6b�ɨ�`eFmD���V�-��̉)�f���lbU�JF	q�O����En⥰1�tǫ2�	KSm��s��:B|�$Ol�9��L
	7�S�Iq�B�v$���	�.��q��O��8�U"�C�1v-12D�d?�o���GX=+����ŦpX%�,�D��=��$�2�	RU��	H>��CJ������Y��H\ip(�����#�K�T��a7���*QX�Z�	7T�ǣ>5Ӏы\PB8�K
�3����OR0*�)Cv�4=a���=���esz�cu�	�A�=�b�<wち<2��ˊ�ZE�D3���}QVF6�:fiY�o��R����z���{���Ō�[&�)��˵��$��b�Od �vSf����.Cd3���3�u�01>��eG7��!�7��=A�15f�����*�}ɀ"��>ĮO�c^���02�Ք�]O4r{)a��?�)tIV�\�
�m��2�
Ǒn��[���0�����`�|g{O���������?�%�>��-��b�9#��M #��1�ЍP6X��o�i�Z��;���ܜ���7�����1���Iz��U�z�-��E�R��p�褂�}�<"�mZ���U�������ւ��IĿ�;+0W��
�K�P��D�\g�7�M���sRa#�&��� rc?#��2^gX�I�g @ￛ�5�zeՈ*�u�L�>��A�*�Z@Z������HI 5B!��*��/ʌf���P�\��y\q��O�9���h����Zf�Z�����e�q�M#�>��C�|����H'50�5L]`�s�&G��,�̩u5�>�&8#T��A?%� V�"�DNX���̰�є�f3p�� k�I������l��A��(+<�7���Nv�{���	�Q�1sr�xA�����6��L2�8bAvO�sdd�E�7��&� �D��,;s<R(��%���{m�m$�xj�����s��##8&<�����`��^�O�i�񎋀v	����#��&[M��L�w������ߕ�}&]�lsK����5��l� �ȩL,O�&��|�eQ���ɜR�EmbuF�[?_jj݄�T-Ц�|�3��	F����[hV%�����D��&�A��V�\�-r��EW�s�؇m�-�g؋�}L��}N��X�*\pé�����ONq>t`vk���B˳��d��Z<��u4��տT�'�wo�ّ�BG���_�w�����11,$9��7:j+fdf�,;I�w\S�5+���W�G��	D5	H�O�$5���x2�VQ��U���a`��g~B�H?ո@s�?O�Ҭ���1 q�SYi�n��b���C[�t��MG��(��ֳC̅UC�8Dyd�B93w�ɉM���Q�Y$T�=[�v��BXl �<�IB}!�!�tWr���xK@�&����H�dV>�ԸF�͆f(�.�[Pa!�|�j�u��1��F�ɸ	55 y>G\ͪM��V��<!3�C�Ǎ�Ò��C�l<��P��T�H��=���?�}�� �N����MP)T�AD`މSOHRmKN�b-��g��ٶ�������7<Ɛu�k.@P�k�D���(����v{s��-ӄ�Y���3��e���C ���1����f�d�E����_k�x_1����|����6ل��o� u����иR�A[�!r��hOe�T�=�=�zo���ءr@�G�>�z�:5 ���KR�d��ue��ԏ�t�̈�]SkV��:n1�~�3`=C�4�$��iT!��M
9��j&�=s�a����y���p�66k�j�#�]�d�(��}��}�FD�^��'H�vw֘��w}7qr��M���;���T=V-��$}���łcT�
'��ύl9��lR-��o��0����y��SCz׎aV�qK���t����I���A^j��i)H	�&�I9�42WI��9 qVY!*9����>�����1G�1b�t>3�E��lU��kB�yT3Ϟ}��4��9������2�v����'�U� ����&�l�!�E��k������>��H�cܚG��V"ڟ��w�yb��x1��GX��&>+���QAqE���X��C>�95č�^b���6��A�?E�r%!]����6���Pʿ5:|�ya�de`"&�\WT���p`�"p�{��A�D��I�L[��'d+lo1I*l�J�3��M�fN�
�?����3�j���Y�ؒ^�'��W��\]������Ͽ������!n�;ؗA��b}_��=�����=9q�	Y��C��ݑ�Y�v3[o,ը��!ak5m��[�|,�����	��"����qaE�b�'#P�Y�q")Y���B���)�em}�P��)�	2u��Q%N�``R8�X?�B�E�������븑�e�q�>l�xh�VP���GE �L�ƝA��"}=��k׈#G3R5ND�O�/.�~,���H��� �*�E5��0�dM����S�����Y���g[�`��A63U:1��8Zj��#F�A��is� �/�`�{'��H�`H΍�ׯ�;�gF24 ݸ_�DZ�4�ȱ�D"H��'�zF�w�d2��g>à��^�_��_�3g����ߓ+�/�j����:��#�hox�q]M��~d�qPS;.��>�|�UM�����T�]�;F�0����dg0��z�*���FmŞ�v�G�s`�Բ�0��
�D���]ge�`NXz�!��m������OK;oʃdo�@k�D���އ�?� ��4�hwb�a�*R��q��ϑ1�f&�g�k�*J0�`�B���@N��<�q;D������ňR%K��}8�a.=dO���bǇ$t�bf�ǅ�N��<���|���U��;vVuoC�{y�=/3��UL؂Th1�7��QՀ�5�H��02 ސ����m���|*�W�6��U�b7r)�L�e[ ��F1䖰��6�����h�8N�V��.���$�\��OZ����*Kl\�1�S��wٮ����7�)�~##�*XC5~#T��lȠ���P�m���r�� ��u "��ޛ_X�9��F���iB5wﮛ��;�:s�}N�����MFpR����������L�p?���~�jX�����`3�4�L����0F{�!?q	�`�Y���&�9 d9v�8���$�3M��?'Z��Ą+�V����?إj̉3q{Í�!$ޗ�^����X�e��=�I�x~]KL���I6_�MIy3�1�d��Nq�� �iR5�`�#wo^���?���<)�bC�pWڕL��W���+r��y��_��?Oei�#���BzHԷ�r;�u<���rdqNz_����z6-�0�8Ӟ�d���E�S6�%��f�e��U���9��OL�go*<�\7*��A%�zm�=�
ȑˤ�����(���d0'F`Ɗ6�����9^�M����Ac�[�J���7}�B0��ì���e��8nN&�$B��^��c`>�|/���Yk4H w��2'�6׷dwk�*����l��b�FoQ7��:^2��^�\��>�/�G�����y-�zG�v� �f����hr�_��/�����R��7貪UM,���(W�������g^xQ����ʅ�W��G�>���w��E�t���hy��}���(�mo0� "�6������H��-��{��h F�v���>92�&1��ҨX�m��+�Z�ɳ!��B�Fm�x��d�IO��D�A{�"t��C@��ٕ��&��4�x))0��$ڌC~w4HY�X�m�^oT(J���tZ`�3n|��R�:��=�f|�ݡu�P��:���q,��*�d�7jV2��	D��W\�[;��9� ���L��R�nS���pnČ�l����$���8t���v�� ��ڕ��ch �:~����P6~������H�Z������<G^���*/^�*�����v����$�ډ]��@xV��|"����:����D& _A�I��(�T*�CJ�!����	�#�����Zs�ߎ�"ŋ���� ��ߏ���ʙ��Q�H��Als�9*b��LQ�d���k�6H`" �E8��U۸�0�f�!C�_<�$���vS�쪼��[�`*�n���߸uG�|�M�u�>��K/P����#�S��}y�9�!PM�MD=/�����]l��C�Vi���26�=�׫�Jօ-c�<���85X�Ǧ*\�X�2C�1�#��0��Q���t�=V(��. w ��.{��=�z�UC�L���I�O��M��ڞ��Ҹ>�N�+y��g(��N^8�c:?��7s�Q��Z�z!���?�r0�A>�����oK<ޖ����V����Hw��ڏ�mW���;�~�&��n�Q�a��P��~֗�7.q���W?'��Y�M["�6=�zp�֝%�2St��EӠ;���:�Q�O����*x0���K��+N;�T@�bG)�>)3ߋ3)n,ʸ$�	M��� Tb���~v?4�>}0����߸b�|1�[(Fb����q�.��P�a�*7��w:?,����t�3ة}NOJd�!#V'T	�X5H�^Wc�Q]4��������ڦǎSCТ��w����޹sTl�!C���1G������Y���*!�F=�zk`$�u�!�4F]�tA���[o��|�����iH}lc����.�>8�����_��Sg(z�,���/���������3��4H��oa�!6~
}��)c;Tk��ya�@�Ϊ7�ig P��"��BN�"����D�Xh��6�M��)(�9}N�8�1������@��5`��T��Z50�p�p����4tXj���9��Ɓ�%yj�k�Xߔ�?8'[[���Dˠ-�O�ZG�9�����~L���!��}:BTX0��^�t�e��Z@)��4�q}u6�x!�B��6�CLr<�Xq�@?B�[�
����ʔ��A#�[vh��z�4+E;m��_�)��/��??��{��n���*+=��C��˿�
�?;3'���N��_������7�W^a ��vgO���?�s~${�\���3�6Q$��ދ*�3�q�����I����=�k�0-������C��*�I�C��IĜ��FX+� �s'�N�8�`E�U{�9g��Ȍ6�:ڀV�uA� ����)~�@��Wz��3�F�̽��d�ux�˵2k߷��}C7h��F H�p�(��$K3v�11�������Ìd�
sh�;	. 	��7�����}���������s��2 GC����Z�^��}�;��s�q&� Z>%�ײ�IҦF)�9VUe��bB1�øn�|�s�qm.�n�� |��Iy�駥���UATN�w�&o�7ߐ3g����{��)(���}r���RV0~��m}����)�Bi֍jƉ��ga;)���k	��ISP�
Bt�pe����G�}�;;X	 *����!�7�6$��3PF�:OH�p_�� �F�U�먣�[�
�~�������p�S2����|�����$)�G�q⾍�y�Ug�~����,����B�L�W����ݳ��1dV@��8��yNIg]��t/���nK�o_���Y�����~>%�����o���M(K��2so������\�uW��6d�\�Gp�P5�Єf�P�[�γ���)��©  m @Lo5�G��d)ύ��� p�G��%v��G�����L�Dl|�Uh8��&�t��2�#��B�l�%�T�p#Qkk�9��ȦU]�q%"�ZOo?G� Nz��X-U�����$�)X0>���Y��M�@6=.a%��O݈'Db�#Ӌ��C��n㿙+&�Bh%��pifӁ��j �'Y���p�ӛ��� ���פ����.n�=� 4&wM��t9�ׯ%6~F�+'O>���L�������}�{g�@gme�U�؄*�M�e�8� �6$�w�Pn޺#�^�(��Saf�`I�{;w��G�}s�㔎+n��+�m��AB�Z�Ź�F&bG[.Bk���K9bp̠w���s�	�C�q����`�1L	a�-Ȥ� �,6v鹱CS�5zp{`�744 ����!AG��J�B=������/�_��A6+�J���𨷌�p����,�m�?c��Z�;�R�Я�~9��A)��2�҈"c���cz,mW\{��xmYr0P54_=��#�xk� Ʋ�mB'�e� H )�5V��ݙZ��%=���k�-VqN�yJ>��/����?���q��S���|X�T >����M���{�]����?��䩧��[3��t���0ᙐ���Mc���#kNG��ł}���~+���݁"��� �&N� o�ii�B�xku5�����0�&Ͱ�QQ� �)�d��b�Tak��E�D�^�%�M+pR��הI�	�!��%�;a��N�ܸ�l�q� i�(���3i��4Q���/H���9��nݒ��y����j�~�	P��[ߖ�w�������3 ]�n�<\�rE����B2����'���ܚ�ӸUe"��(��	�������,3�w�g/��������!y���ѡ�Z��D\^YeE�Ur}&�=�l��J�V�k_8�^*�k��:>�G`���ӎ�w�������Sr��UY҃]�Yǁr����. �$L�85�0�̘L{���y�krz$�4�nV������������l����E�	&5��n��n��[u$���-��´<�䃲w�nJ:�.,ʭ{s�w�V�x𔄗.�{̓f��㗥)��9��)w�~�gӈ���zNLK���ʱpz��D+�����$��Sm�gI9@���F�}�H�I?��#���C3SM,5_�b�rRL��,�E��u�,�*@��<涁�je]��2;sW�EzXl�X����|R0+�<�e��S��и��ګ�~����)	��G�L	��2�׍�L�U;�8�f-�_g3����N�S�����ZV�޾nE�yi#�.�=%G4T���rZ��t�s�{r�)�Nʁ���¥++G��M�%�;o�SW�����,g<��255�C~5�V4{mC5}c��Z$��Mm��f�$ē)#���;���}A���7�SÔ&n�t[*�A[}��Nm�Ϡ�QV ���v���xT���K8�c�|�r��#��0���W�i/>	Z<��{�0����Gc|:6�Lܓm�aDr��]9}����3� ��
����:�\�$�"v&fiZ����X���!3/ߴ����b�4;�Qĭ��KAK^�z����ْʊ%y)�&���xT��˴��v��t�t����\7�<ߺ)���D�|�Lc�y)|^��w�}p麜~�y��_��oU��]{Ȅ��˯Ƚ�9]�W�]��ݓT~��r��-���`pB��Sw����c���+EL�xD���@��8��#�a��"b����TG�����eߌzF1�QL~�-d܇�*��f�� ][nttD���c�a�s��e9���&47�ߣ{���h�\�tI~�ӟKM�}5�&� E��X�����Ϧ��5؜'��6�}6r�$>$[�H�%��6s�ȩ�"�����qB�� E[�
9qPŞ[Z����,���'����2��L��&���f�W҃���\Z��g ��.��1*��y�LMOK���C��RؔC
N:��O=�Cvim�E��vu��z�ͪ@6*���8��'q]߆&�9j@)`�����Qd��x@��w{Tʞ�se�������I���D��].�3QdSJ~Ԋ��`�2l� �OBzߤ͈V��]٦�C*��P�Ό�^��YB�7Ҏ��6�!��\����} �v������<tl?���Yc�F���M��O��.^ �����V�ڛgei�,��_�3�O�N��솮��>����Y��rVUr��s��!����"�?���[i{�����أ�M#K,�9�d*���hP�4�*��\��"�K�2;uK��iVR�~�"ʤf���y�$ۨdZ�n�mSY���ƺ������Q͈���êNҲ����;�q��u�&��1�n-V�W��8�&p�g+���b��>�b9yB�<z��Q=���ώM�"9��'ΐ=TZܪ2�a�a �����8|pБ�!�z�RS������]lY,-.Jp�qN��+�d
�D��M%�~d���ЬLO�VR�>�ć�*ٮ	�Y��@UN��z����HhH�%�,�ĺ�W��Ald1 �̲���|� 2��Vb&�C�}>nw�E�c�o<'N/Y�UPI��$�YU�$xS���n���o�>�|�! 5�}�j�&+��$�dj�c�L^�jEfEۮ�83���H&9)D9���
`�/�.kЂ�ZVAe(O<z\v+������Cg�tm�9�W&!��Ո��V�	��Ŝ���R�"��Ǣm䐡��L-����[�v)T�.%L�����3 ��^)ip���ǖ&�����!.,.˝�)��.Y^[���%���zJ��7r��yYY+����w�#���N ͪ#a�s�r�e%�H�v���س�G���~8S5�tlY\%�V��E�!&ɽ�6�Į]��_���y�+��L��3����~[����TK��?�r��!
�p~��Ʒ7_{ݞ�S�{V�.�X�VbY���H�ݛ����]-P��U�����1�&1�Z�b=  �Z��l�I�� ���^�K"ő�
 ��(	�0BCN�|X���/˽{�r��wM�:
Υ����ۖJ5��H0����խ`� �K�z-99����I�Sg[J�:e��M&'�dzn����}�2�I��S�Q���/� �{�����y<�6٫1t��W�' ����ϫ��<�M�x��=���Y� �gɦ���������<�\+o���=�r��M���g#|�H4R>L�t����Wa�̷
+����o�"��eDA��H��*}�I��8!u��%?�����Ji;��bE�u(�wKcy]�LMd����Zڏ?��<���������Sr��EV`��g�W��ª�I�.p� ޔ���T,���c.t@ϧL���=O~ˏ�����d,���Ff�G��94�����ܻ}E�����2=t2��5Xt�w��#�IP�����s�'o�=�M� j���LoWd@AA��n�`N\ �@'�uBhIC��
M��T�V�'r��Q�&r�����t;0m���%@<!/l����qVE>�9wV�3��߅���c�kfyDV�7���;$�������r�(+
P�o����կ�$��k�J���x��M���ʣ�>��g����{�� r�)W�%;B\:c���!��5��k�E��R���6[7&�p�l(����	}a����s)mlR�~uu�T�tK��@�!�C�;c1�P
X��H�K���FuG���M²[]�w��Ɇm�cGjtSZxN�r�b�#8L^��DN�$�"$�Y�����n����V���[r��a��}�u�~��1,ϯ�?ܣ��S�˨�U(Y��&�WS���"B�L"��%4ۀ�O������rQJke~�L���@߈;rBfeii�cø&�+P��s�(�k����[�鹩LZž;&��1E'��H��-U��~ZB�Y�fڐ
���ܙl��ipp��ahl\޿��S&��435��R@\��o@A��������`s]�4�JI������}��B��:g���3�����?��W�ڝ�7�%�[[�� ����,:R�����~V^{�%��w�C�O}�Sr��Aуሮ�����?�>��p������g&�z ���yN6ћ��Q��u�8�=q�k[�5{�Q�Y[�	�����i�a�3x�u�����˫� ?��;�C�#�gĬH�ᥙ��9�<���ɉ����P�2EN	���	q���rNr)�(6r,��\GGN�?�����	��Ɗ�}��S��tud%�k�|�G<&G�;!/��E�}�A�W^zI��*������*@�T%����"�/������Uj�`b)I7c�l[|7��K}Є�~s��n����Q�y��������C���G\5�M�M�`.�ܴ�Ȣ�5~rJ�}	�XQ�
��!i]����OߔZy]A�Ga�Ύ���?���T��;��G�� tx8�
Vl�o��#G���@/+��:A�yo
����,����ے���<,<J�7��s\��y$�%�t��^`"��bx��y����c*ACs�1�����i�VED5 �������R\�W��M3���NٻgRƆ�9UQ�Z��δ�����[3����5�Cj�k���%�s@:�:���x(?���V�)aM&���X�4GT���)r��0j�8P�r�ۺ���A�I�f��E]3h,|TNg�f$���SD�k.^�(��� B��/nU�l���n�����V��5�)���~ϒ�-/�BıP�/~��������,������i�v$M"]dx�`2 @��`	 ��L����A�z�v*p� ��ȶ�6��t�M�kye��q�Xdg=u�W	GL�8�@��,r�ꄛ���šE�Е������;+�]P�m��� ���R͌�t�|�n��ȧ�
���[�ȑ���Sgdfv�َ\�l�����[j^n��د��۹ɱ�s^�r58��A�!N�JcK75�{����G6׊�<q��k|����9�b"���ʺ��3Fv�L
1EC�徍�k]VY4m��1u�q�&��$sC1A��
��]"�m8br]�� ��=�|&�k�v���P1�k�X*������� �����̌<���
�_�����F�z�t&~�ecv��:� �u�V���5qE�V��ȴ^sڠ�,��w��Ā��q��k �R �U�P�a��/�݃�:7=#����90�������d���jԜ��Rn�P���K� {�n4۲u�F�m�'v��3��X7j��-IH�Q�͔����:	X�;�*����!N��k �xλ��a��˗��<y��<�����׾�5�����0�c�<nkFV���S�FE�́�q�]���=��R\]��a��,֤������ItP�v;�dh`��.�(�B�H� �M��O����������#C��6)Ñ^~�2N�wtɦ��S�H�MKiۆ	�\6��ȭB���v�����}�@�N<@q��]l+�����))�-q=A�b`H�C���n��7K �@�jKf���*J�p��}�z������
�G�H�=���������_^]!?�h�"�[�WML��z��V�
�Z���Y924*�[r�<��ҹL?�1i��:����������E��s�c��)�E�W!�� �=@��n,/ȭ[W���L�i��kX�9�V�<��#��D��K_\��N>(=���O��@��j��Ս�.�9]�	�#����T���恘��
�hǏ�]Z�8~�{8�B�**�8\���Ϗ��Q2���c��Js�4l����ptCt�@���$��鍸�o�h%���rV��~q��@wW3�o����/_��]���(u���JZ,��Y&B&*F�Ǹ�6�����4�!4pr��不�N@		����C�n
�f	��mÑҌ�@Fs�9P�����M.�㲡q���^,���dy'X4ޏ�r�h?r~I���?����,���'�f��6AN(�@��w�ɳ�>++���k�����vc._f��i@H�}��TtS�~��E����h���#tʣ����#�obhB���d~fQ�|�)y���2?��A{��	[�2��D��0K�xb�#�'�x
��~G=��D��{ZF1��F[6őp�I��m�9M�h��n�[��1esm��B菏��˱�˂�iL��M066"��������������׮���'��3?;-���&�Rn\�*����xv����o����ˎ���.i�&�Qb�W��a��=Z�X� ���D�!��O��^��\�n�|�z����/�#G�ʊ����(w���*li6YUuWv���Bs�ִ�Xg�1���X�[�n�5l�WZ���a��?2<���/�&���[� @e�ĉ�/�>�X����?�� ��,ȉ�����r�]��yg\�ݼ!�[U�j�x���Ԑe+1\���Ž�g�27�v*��eKyZ��Ҳ��)�x隴�^�{�����uV51���;o�!+���:���<W&F��o$Pk���`�?~B���:$c4��h���o*c��&�4�b ,�[��ȥ�
]$��|�Wd��n�x^CRz���IQ�;�/KiiJ�]�-��ʼ�*Н���&8;�fњ- (��q C�]<'��>���We�P�/��W���=��?`z4,^�~�9	�ɝ+/h�0�
K������ժsR��3��ۂ�Z��qE-����;�L��XH�`E�[�S�Bm3�O��0�0��G>>v3�Mxq&k�a���&͋�c#�ܺy��XQg��з�40der���uu�}��T�,/w�re9tx�������.����4��;;k2����Ϛ��]���Ko1C{�y(��� ��57^����0wT,�h*(F�ā�ʊ��PF_2�؍�d�m�i}���aN�l`�h[Ȓ׬\��ZgFt��)=S�hTK�lx2h� Ѓx��ɬ�����n�,�|�,/�_�$�
��a�/ ʠ�n��8p	�JF�N���!���;����_�!h t�!�#���A��f����P���d��vr��}�9�Q\2�±#��w�|��)`��+M	��m8�:-���]�vy��
"��{���wϝe˃#����%Yj,���C�ZY�3��2�V�@�E��4Hu �I���FY��-Ք��H�I��?�g�*˕�פopHҥ�x
d�9e����<���R��a-��i�,�1�g����l��gA�OX�g(CK `uȺP%�Ҁ��9��������Б��/��s��{G>�tQ}����?�'�?IB��ĸ���/�==z{��r��_due��d����G^�ի5���2�P�L�B#c��Q�� �q������Ӑ���+^E��S5n8?���Vl88D)�ID�
������GkQ�����\cV��"�g����g�ׂs8~�^,����xb��0r�D�v�nE;2}+��7b| �ۓ��ܬ����zC�:*�.����g�zhb��[��u�&�<���4x㍷h��ЩG�Q����r߱c����w��7��P��5'����,*I��HJ��GU%���ho���v)�(m.I�ƈ��v6�y�gu1K�E���5�o' �@j�S���G�!�2Yp���&W���!\��feg�ң��|녊%K�q����� f��á)��z�'L��_�t��ВD0��hJ"�]#lx[��3h��*�(-ωlmH"�3���jyKfu]�:��T1G{T��n\����b��K�sQ�G����K2=7ˊ����t5��#�'%<C�r��my���$�"8C�ׯy�}	-�m���X�7�Ѳ�Z\;����ѸP��#�z�H���Ƌ����H�o7�_�Ձ�LY����m��U�wC-�a��O>��6�� %`����p�9~T&�LȌp���PIO��z�@0�]z�;�S��B15O�OB0�؎�� �{�0v�Q��7k��l̐B5<'�8E:&t�����F���Z�(���R��#�*�Hy�+M��,`��)�Q٧�cۇ��"�� 3�F�
��GP�|<*	8�L�(`���) �M߽��2!���2G凪��Y��k`���\��aX�UX�����c��6o:cc�j`��S ukv#l���C@�F�~�#�K`3"bq�I.����Ob��UVL�ޙ�e�r�j1AW^�9	�}oc�귤�"�a�w��7'�����Z!��x����`�:!_�����'O<yJ^x�G���H_���
[`�TN��<{�Q��$�RCʛ�re��?������J�_��������?�]��&?x�yfs Q��#��g�a�����
��P��������*��җ5(�p-E~��"^o��31 >���g��G;#��Ʒ���6۩�d����↹<�E����s���	�!��覐�������Y�����_���1U��˿��ڙӏ��r��=�|��f��s/Y�cōk i������aʰ�j��(���Q��H�3���6�k�E����0�C&��D&��%����d�@_�T��޻�{�����yP `?����矓���g�E��t����;�qr������J��HP,n{���sF(j �h4�9�q�!�W�����Ekw�P�Ⱦ_������Y��q_�C�L������5R֘E�p����"j��:%1S�ȑ*�K�YxMc�*��cGIW����xu����gO������=|D^��/edh���"��'�
n�~Cԩ��V�Oh��聓��E�����k���c>ER�JC�*鸶��v�2{.	J���絴s�f|&�h68�D�;���);abxP��Z��[cT���
�i]O
����|z�A��vU���{hP�J29��k����QL:�M���!YE�4;3��eSF���(��#66����0�j�	e&(L�pT�~��qɵn�1O��j�?8�`⊶ke�,���H�����
T<���+C�O�ۤ��A�/��C6��5jaj6�bڔ��;���9f֎��������ܧ�׹wޣt0f�7�bTQ�߿r�UY&�hlIowJz;�䁣4��͒"�D^jwVH�9��j���uۍi�{
���z�uҙ|�~��@��d���TiJ�#-�S�Hs��bb�d�����|�s��#�>,�?/7�^�I��Q�fc=]�4\^\`@dX��d#�}[�m�@Jd��}���z���.�ۂ�ҭ��SOiF��j@8.�߽�Mo,�'���{� ��w� �ZZ��)4M��tb\Y3ľ�N������ �����PyU��f���mY|�b�&��
��Y��{TU��%�qx5�C��b
�dX��<��Vr��ޑ#��"�{�)��TJ�e( �D�x~��\�}�)��[7��ڲ��G?�/>�y�ʗ~_���_�,����H6���]�}��؞�z�m�ނ��}���IU�!z��Wg��/��s�}�Bi��ޏH�|��'eh�Ov������C�dF� ��߽�D���%͜��f,k�	0.�c���
�( 3�������������U���P��?��6���Ko�,(�B�CelS�T�Y@���7�#���w�@��G3�������_	�q�szA��C7+��� o��J"���8$���L<����5@�HZ��o��ȄDk��b�1�br%�5/(1������k]TP��2� �+k�z�U����g?��dǆH������DV5�J��ǥX-sD-ׅ�e]cf�*̌m�*������D��+�7�l�I�i0�M(��O3Fs#�*JC�$b$W�I�Ж�}�^��#� ���@�x�<ï����q}&P��x��~a�]Lj���mt�e;U	�Й�2j�w H����pD����L�\��8q��Myd�����\�~��ޮ�>)�Ҧ ��n|��+b~n ���R>ȳ�==�^��ʺ�IVSSm<<��t�B�@���oԈ��|ghm�؁�*X>﹩������?&���I	�}�yS|�D?�?;�LZ_��Z�\)oS��?�P�NS%�tm�a}�bjh���dc;�������ɼ�$ }x�a���F�Ǐ������X^�ǔ�(:�8l{vM(P���A�1U���;�	
��ӹ!�N:�s�nGf��$�^cн�̝��z4��ߥ��z��h���.�eV� �L�GfӨRY�\\�Tʁ��a9� =G���0nPٷg�,�-Ja� ���2>1����օ=><J���Ѐ1����t��<��](��7�u�PdJs27�����C�K��4*��K%�&yMd�����;�b� ��,x�cC�5�YX�/���8�х���h'F_���t�Lk���Rw��H�� AH�L:Q�wξˬ��Sr�gU�#Th���2�?,<t�+7nޖ�zo@��T����\�������w`p �����ƶ��t� puC�C3X���%W�J7a��`%���v�)�P�E�j��[���4��c<�L�ۮ�i�o	�n����������&B�Y��g��vj"�Ȧ]��\׎2��7��CJR�;𨗡� �D��u��R9�^�#l�W���48~��OɓO~B�L�W�K�u�2��o޸'���kr��a9t���ާ�<IB+ʮ��lF��5'wn���Ƀ���$ǎ��k7n����!��F=
�q@"("�k���2hܹ~S.\�@3��;�����(�}��.��+���^}EN�~T����<x���>-���7emiY�����D�}���¬ �\��`�h+��Y�C/�7�Pl/$�M)��Q��	�V>��"�L��S�~2���D�xE0���Q��+^p��c�a�a�\N/��ǖ��ƺ�0��Z��)tzF�nHic��FA�� @��iDu�K7��~�ߑ�~�iФi����;�����(���<�'���c�E���E=8YU�d���k�V%%^�Z��5m"ݮ=�u����ք����{M>E��^�)���'��$ �Fh�ͮ��z⬋g#��q��5�od-':I+��mpt�{{U����)��y]k�\�8��qi�"��8!�]�n�qzh��885w���
45�zINA
F|�hu�@?�#iR��|Gs����"�J� �o17e/�����{���o�` ]�+����W	���Ŕ1=��KA՘�c�JQ6DȮ��eB��F��o�I���zд��Ѩ�N��*&�4��ir=?;˪74h��G���;>
�!���Vo���8�&�O����ba^�WM���$�׀*P!!����a\J�G�����M��ekM#AxQ�;&�D_�VI;˘-��e>���o�JA-P��(����yv2\�!��~wo�<��)9w�])胆����,-,I�KI��Lv�n�)N���#�ڦta���kֳj.���j���X�����	��g�'s�P֣��Vyȉ�_-�D͌
5�P��C�'+CÒk����}gJ~����ȣ�ˑ��Q�@	-�v�<+k���O_�+�nХ3y������V�Q����$)�����!�#�� �\�΀
]�d&ߜ��ؽ{�,���2� 8+x˴��edp�zP�eR����0{�K�32�0�YX'�a�1�=�vk Ue��6N��M�����e��# ��t!�ql�1�Y2v,Θ�)+U��I�=�NL24�J��b�������C��%\���0p����OP�VC�jIZ���*�my���������̓�˧?�i����_ʅޓsgߐ��zU^}�mfs���#�zIA��.1x��ʟ����������ʑ��/�:���M&?@z�f�Y]p"�f��U,(�/�Z�w����	��<����fC��WVeM�{S�*0��>-���c��@�ݻ��忖�qfS���U����V��_����6�	C�,-���3���N³�%8�Mf"���s���ŢY�Ԅv  鞃J(�(��ۮU�� �W�{ ɼ-�&����s�j���g���L��we�"0�SaqA�������,�Z� 8����+�'��~_{�_�����ܾ}�5�C{��Ҝ�G�}��T� ������M'�8�z.��Dhj�������Z���qyIN	��U�bv̵lX��>�S���Y�X�D�� nl�_�aY��'�͡�����wdX�P�.y"�'�g�.�0t�~j����-}�5Si�*ھ�fzz��Ĥ$�B���� �׽D<蛃��%_�yV�.�D��ԼW&�g,��E2Oϳ�^P���z�?И�=]F�D�k��.~�BG^64��:H�<r\�}�^(��iz-Z�$٢�( Z/������ n�}ݸqCAN?�2Ȭ5��p 6�1S���!Q�DB<5� f�*�
T0�U����6E�pJ�s�&Y)�
-��o�&�j���iłS�Ӆ����|�@%r3q1GE\9�}�8!4�2r�1�k�>Fև�W��.�<{��2��.��5��]X�������<�G>"��\��Ӳ���1���n�]]=�A���R�Nh6�,��M�`� \$�ᑳ�VʊD%�}�U�*[����@���^[
q.U���KTP��DS2v´������?yQ���<v�a�������!��?��/���=E�r����)$�Y5d9u!���l"��ˊ~��?yA�~����(�����2��k7t�5�����oQ3���L�@JL4L���+1c/ܓ͵%)�{�������ԩ{�
��`�^� ���أcCzh�1jlp�a�ܾW!�U��h���93��9g�%��9u0{�$�r̓��
�9�[���Z,P�qy<����$D��p�
�A 	��jFuZ|-KY����4�_���\V0x��Iy�SO��Ç�����_�;y��| �u��u�R�=��]��|�slca��k��m�{o�#��=N �'�:�H�e��0p�D��O�9Ҿ[��s�sl��(m�<��j,Ղ䉲22�l*����4)�D�I<����.j�DѦ��*5�D����"��Ʉ�n��J^�0�9��9�L4U-C�¡�_�@$'c"��c����*���ə	}Li� l�0 p(
�ag��h_�	F��bw渕�VE59�w���M�vE�A>�J�[o���1׆�l�&���w�k�\��m�L���4��!��OPmN%��f紓���G�r�O�#_��(gS�VܶL���E7���F�̶J��=t�߶��3r�Z)�gKkk�U@��K2�	��P[�gӚt�A��_�UMچ�'e��%9pR�8����'���+��N��B�(����]&�����~o�A��<�,����Y������w&�"�ʯӰq�;�`Q�����G�
`�F���smI�u��ǀ_��˨̷�ۤb��>M86�n���D ������8S�����|���M�ڐ�7�>�D��U�5M^1���e�AC< ��c�X�Sg[����ȕ�Wh
�U�R�S���T{��t�"�FŸ}d��Ꭹ4Ӓq�;>g��Z�H�gZ?^��R�d@!����cA���.�ϑ�s�M�@���3/{F���{נ,.���윱����F�엿��L�ݥ�~�6%���_"]s�K
zn��Y�ϯTdv�$o�wI��V��k�	���P�J�,����"z�E+�q�U9�5N��c�7Q3�s�e�ܨ^�*�"녀�[�U?C�󐍃`���Lξ}��Lu���'����Ս{���g�vW64�.)j^^��ӆ.H�*�}_֍���l�vN1���U+�����w(�maWm�3�d�~?���lWȚ_����n��GzL�V����S�� df]���
'c40T4�CtF�ﹹ��(}yѤ�1v���/J�#l"�� E�`��C&2']d�=NՔ��&�\�Oc�ʤ�d7�gn��9 ٺW��+�l�m)�o��%D�9�fK(�»)I��I���U�/�"�ο'G$p۽�਄����[�.��۵kRAe]���K޿pQVVכ�[�Z�!��e�l�8��1��Ս��u]�mM^�DE�o��?�[c��!�J����XD&�������v��ͨ�I����^D���-��ޓ\��@$�-��ظ��ϭz�J3i#Fc�����D��aU7jg�x����+ŕޛ'�~l���K���g�tͅ���i
&'�z����G��32u�&	� �Ȗ�E��.EWw��u���@�<t�~����k�k�Gsx/E=p�DP��	"��(95 \��>��U��]�J�����L��Z/���@g���z��zM`d/[L����
��\��N�7��_�e��&���Z�w|��O>Z{�K6�'gS]7!��h��diG��l�`���'��#�7�K�ݾˑ۱ɽ�2���������ʍ��|�чe���R����w�>:����ʦ&pUM ο�8�c���&M�.��mK���ԁJ7�k������Q9��T`X
"|��Fa9��`�),�l���
�ҩ���K��>�WJu���p1����WϪM3餂m*��$�r���<���d�������A��o�$k4��/)H�=�wrB��W���K�b m�)�é��uA�qhTcR���Z��%ET޵�e���C��<k��GV�(�g�mC~ۏ�����z8�־�\�Y�l��0j��@"Ҡ|@˱C{�ч���}��AhpP�������du�:93TL6/\`Y�þ�~iנ��d����*��
T�6��Ԣt��џ��M40�ڨת<����6d�� q��^-���t-[�g�6�;O1i�+���v
z
����)m��Ͼ��U�c4�^'[%�Dn+8��������ƞG�U��|F��+r�*Ƿsm��I2��0'x��(���)$��Vz�r�?[#��ѿg��<J�
�:�)��"W��әNc�
���y%y}� �� .t��e�J��݈�,ϳٸ3Hͩ����xf�涸�X�*��*H��GōDr��?X���ȵܘ����B�2���MT�`��<�Nt���9���iB�E���̶�85.��i�g6j����6Vm�D��
�^�#Wo�e�D��: )>A84q8@�R�BY6�e��{=>:N�S\3ڤ���
�&r 4����	�ξ}�R�x�68��yB:�I�\�K����ܹ�<����/�<�}wl>,�>�����/��ԔY��#�N��ZCn�;JpD�Ƕ9����)w�A��3m�xt�¼�Fk�����=VcO"�� )?aE���.�ˮ={�����}p��m9{�N��Aݪa�w��!��н��XV`�,�3SԎ��s||��7�М����!L2��Uĵ��tG�"�8�5�x 9���&�З����jɇ	������&w�}���ɯc����|M�D<V�vVO�0�gm��x���8c��T���#mI��u�i�߂V1Y�LIJ�J\��h�ݼ7���ƤM��tG�l�!I��CpeV�~EbL$�wI"�!Q%����(�k���{����|/��J��r{f���2W��BK��pf��F�7蟤�^t-��I��|Kn�e/����B�J�ɠ��W��'��R�����LѠ4�nHb�\���9oj�	n�����S�˴��A�����Jii���/^}]�%���S�U*������|�1�ҭ���{�4�������V�@C�˶�	٣�^NH�J�*�/���Sq �F�LrB�iY(�����u�%�+Piӧ����"�X��k�Ɣ�,�80��6�46�\!2ܷ{���ܲ�N�e@�;3w	F^~�ey��We@��	E�{&�P *�ʲ��R��i��͒�@�j<c�	A'����M��!F|�g�+zN�n��w���y.��w��)n��3�gy�n�0�%ܸq�S5}��j�3T��>6Ҫ�Wܣ�f$k�#����G�nn�b44��g�X�!V�*�h5$��fZ��SO_?�bi�����\@ �@�����2��-wo�$���Xf�ޕ�ʉ��]#T�䴐o�"�6��b�&�'Fy �s�]y��[�])0a����P2`��@*e�*� �q�:��p;���pA���\`�Z��+�h�����랙����2�X�(g�m��43]�ք�!��%t؜�X�������k�Y�;��z��\-�Ӑ���	ΰ��VCp�sF&hfk6��m�"QIz�6{P�ٷG�eV��M<7eV3���I��|v��x�h�\�qG���F$3K�%�����_��WTY�v�2�d&���?H)��#��3Y�q��-�4�E�Q�Q|L��V'�$��8��Ăqy��	%-p�0��6&�'\��%2�`�U�(Vau�"񈱫�%�u�~������ܸ~�.��@��Dq�ɺ������:�ö�e���m��(t�Bm�]N>� ��.\��_ƙB��G_:�'y�$
}��C^�l(��!p2��!�)�D�0r��&�(���j�;���66\��F�cr�9n۔�G���X�J�lh�_ܳ�{G�ɴ�= {�RX�x�u r�$�OQM��@dMJĝ.�\�;d�\����U�qwF��\�v[�6+�:u��E�]�$�?4J�&�XCs
B������֞���1� m�$yi�V�R�=� �<�B�'	wd�Q�G��լ.���d��w����\>�� Tr�I�]QS�0��/˿#��#���W�	�U�̈́�=�eQ�z����;"��e��H�k���Ɏ �� �m��^�ݑ�ME{��}��m���a��)UzVt�W��`�&=CVi����`��x�ۦ�qI�Z@v.&(��s���N0��W@aKg��ߚP���i�Dr[3���|�Ϭ
�V"&�?H�����1Q�Ń�#���4z�`''7��=�����?t����8y�!r��p=,ʕ�D�J:&��ȍpY� ���P���O�6��C��	�Кh�Hܲ�ܹ�r&��!�U�hצ�,+��$A"��AK�LH���}�T����m��5+�)zf�$|��V�7�J��5A���64��%��΍�a
�Cߐ5�?�q �[_�^��erlXF�dld@:sY�W�����\ܑ�G�����|G�"Mqw@�����љv�E"��4_kttP~���<J�4!\x�����8��6!en�[��p��h�&��6�+����P�ˌȕ��ٖ3n����Mx/𧩡���I��Rآ7P�feh��A\��������k���w^P� �^��B,�x4f���c{N�hBg&���Gn>7����?�	uO$�&A�-�<�Nݑ_��%�
"�x� ����uF3�P�:n�.H
E����Y}�������е���X]���}�� ����I����	��0��@�XD�e�*��#�����xqv�bT�����!�AӁDV��AZ��)9y�A�믿.��Lj0m�B�1�c{;��E*� $�H�ɐSn*���4�>���Qx�Q������A�ʻ����eI��%� �M@�Žf�#��G[|�4I~�;�!ny�ﲣM�~��~�H�[Zu�w�����s �kN7�,��˰�/N��Б8	z�D����*$�A�hܦ��m("�O.�l��Ҫ��������V(U����kV���_`<�(�$�7����NO��h���]A���4+m����F�&�H�$FtS�v�u!;Gf|��z��9@?��gk�����yP�ầ�>$�Q��b`9eURN����	�؃���Er)b�Nf8�0���|J&�f�s��y}�4����m�8���;����|[�a��s}��2�gR޿qC奄���TW7�|Gv�������WD-%����<�k	;�~���qV�4�7�
+���d6�|~	�&������
��FL���gGg���ݓ;���L�����+D�P]M��Y,HBz�V���Ѐ��P�*V��wH�x�	y��7�����Wd;J�Z��ѫ��]���$%�6�?[�T�'p�K��`2ץՀd:���P^c��L����& �|�>l�`� G�:;uS�%�fք1f]�5�4��a�̯����k�:�&�}z�d-(#S���W�y�R $�	ˊ<:���?�6@�dzf����e�TdV��NOw���=�푙�[�o�$�QGFM3bϾ�f_���\�LD�Q�	"�(�@��;z�ݼ���w8��'��o�5	� Uؤ��N .�J4yT�M'��0��٨;S1|�s.��P��3?��Z�d�7��R�����k��F��!s^*0�A��1��V����Ir��T�S�f�:�%\dl�����a�Sω��#��0�p�=5\�s�%[��Kd� �!�O����ޞ'h�L2R���$ѯ�x�6JȮ��V�:cB���k��$Gi[�w��u�d0��ZSL*,P�)f�#)x��:jڪP��)��Q�{�(W%�w��hz誛�F;8,�e[C�֊Ƅ�&���P>��O���|��`�J|��#Ԙ�����_d5� ���k	�Xv;�~$�Cؐc��^�\�(�
����拐Ƈ�2��Z)L�5��J;���fI���b�oX�Y�%�"h���N<Y9�Z��`�����=a��w���Qiωb� ��Zښ��"�ɞdy��Kq�9�D�ڪ	���=|�1y��y��c�#o�=jok��ɚ����.ט;d�8�`���*XV���b��IQ�AU�Fo�SF;��ɠ��L*��f�-��ۏ��A�����]NH��C�P�Ƴ�XK��� g���x��><� ����^A���$��3��u�4��G0���p	oT�P)ɸ�ʄ"�(5��L��y�ے��> #(KP���3*�pK�e<����kH�֝Y ��u���ݾ͊�f�z������IW��mIz���+D��1�ó�n�c���B�_�xq �{z�YK��,d&|�w�D����D|Ȱ0椮c�זĵ�,��\;μ
بOi�mo�|trRa������
,���v˖�@/�e&��]tYXZ�U=�6��Yt�]�����rU�u��f@����{ϠD�<�2�m��П��En:~�j���cf�iÿQ9�?Pv��L�(,�A�'8�K�Y��&�M]���<ƪ�&� ��`��9p%N��)����-"�z��2����t��*0�	����.���jGwG^����s��i�59��u���c��8���4bK1X�i��q���K��!͂ήvY��F,��DaNH���pό��d��=W/���+]nI�8ʌ���l( �r�Z<p���`Y��U#�ݦP�����-�,�2��h6B�����^_�a�d̘邬�s~TQ�6��U����#�Y�'Cn�	���|�� $^}>8|0&��$9*[�t��%��&�6��ŹU��sT.m���us�U��8�لU�
s{��x/p;&�XV���"�s�:h�;�<�U��B����>'112¹s��!�f�&V�9$�ȵ�W�M��6��(ǒ#b]\�G�;*�>vJ�߼.o)0ۂ��m�+$�J�M���ۀ(J�XK���ch��	1�m]K���7xkm��������B���e�kk���m���{ǲ�<��ĕ=W-�ǈ[�4����X�"7�>����K�۷G�Yq�E��\�$�v��`0�lr�z; ��mA�M.A���ԈUg8گ �ڐ���<q�1����WmbN_
IZ��FC�DR������ ��0_���9r�& ��^��q���I3�-l����i8�>�6,�q�Zպ�u߼��	�h��6������b~`N_L�G�$	�X��:� NA@������R�;3Ѷ�r��,���\� g=�5G���8&p�w1�mH���-�����=��rW�asᮾ�$��jULá��ʷl)�Z�@�WN�Ϲk�dK�#h^G����H��n�蘔4���_���sq)�En�ՁdI��4Ō�c�dq� �_*
�$$��>>V��%��N�ܰ�/�ǖ���1Ј�"��A�P]��_�y)n�p�K[�ҝ흒��ś/����"AY7 �&�n\�H�gߖ���}@���fL�d9�R8 ��e�,�Sw=�(0�VPX�I���
 >Q��ck�z�����q@8hX�%؈߻^#g�qy�D�����P"�J���m����2��#�=���lNQ%�� {kfn��V�?��I�M&�!޼qMz�sQ`r��
��t*�@0�䧞`E�1W�'��>��]�y��w��	�J���)��gϤ��_�%��㟱Bd�vH�� ���|O��*B����T���S�Q�&Xa�7e�*� nzm�0��GW�M���^#f�K3��N��]r�}����ʺ��"�������lj
�37LB��g��A;ƍ9&���V���H��G2q� $#ݚ1��nG��U͔�9B���}{vˉ��jv��-@�I=w�]Y\^!��ς��1oh��_J�%���0�Z�W��T�YK�!%�R�I���,���Ƞƭp&��I�C%9��Zsx�KD@��;�������$[��sV�<qZ?Ir�����/�9�{�yk ���ѧos  �!�����:+*h�@��\#}k�w��]k��h<�z(�?=u��DX��-ͳ"����6ߑ�ER� ���@�$!�Q-�BI8.����� �2��}4�9{q�3�Y	�<Wܴ�^�蚶dv�[��9'� Α��d��-V	������� ��y�
��=���b{��kW.��G�g�
*b\�5fՏ�ʆ]W��VLE?W�}P_Za�ئ�_�^K�̠�qEq<A��t�*�rR�P2m\N�;ǳ�ҽp��=N@��(a�ވ��Y�Z9 �Ve6�?$`��ֈ8��Gđ^?G�*?�~CU�8ݽ�R6)W��j8�R���$���#&����P�9���Q�n��蒍�i�m�k��3t�S�;�{��gi�Vf��/`"IA��L�Ф��������OH[�O�7���4�ɳ�KFpn��7�}w%<&������鞠{8���#V��������'��zUu#��8*1�)D��?&���u+���#P)W���Ү��{yk[3� �}]|��j^N>p\._���J^�f2��k�}�iyY���krXF��5�TX�b���h)^�NG����V%	Rl��M'����m�Ul��ƵH�������`g����I�L�
 ][:�T�4_�P0�h��w<�ja@,#����w�`���2O����D��=1I�¥�i�@��"��yDz�d��k��7m�VUl�A\��k�^=3Z�d�Ǐ�'��J��/IgG/�&�#�£�%x|�P�{B�K&ZSV�je�6��	qul��FQ�0������1�̋5!'Vd �����z��?v�BJS��p}>|P�����>�����*�!��d����6�>LR��փeII��H�G��AT�4&�$t=���C�g��<�B�섦f�m9�7V����k$���-iO�<�`6�]��'hC�Z)�}�: ����$�c���^�����v1W����%V�m�n�q,��!7�CW52΄&��+�� �A<��%Z� rیʑQ�	V���駟&��ܹs���fR�Q(�4�{h�`�-��\��P�� �ef��S�R�@*�T����$$.�7�^��� �������JNR�F��v��E���\�ud<S��*l-�k\q1w�f�%&��� yN�-���iy�㊯;�Hb�y���M��\�=1r�u>��9 �@� ��5�q6!�y5a�}�k-J����)�s�v3���Eh�X��8I�a�
3>>">��j�m�M��팙H@��َĽ׵��$��P��i�j�@����U��RF��<׍�Wo8�%���iL@�i)p=B+��5S�g��P�EF2	�5�V@��
�*��Q��Z#�V���� 0�S��Q'�X�%I+�tRϴjC�Mһ�H��P ���/�K3R.�)� X�#c��C6�')�3����3��q��K"�!ŭH�ۛ�Рe���V��֕4[����uEVBE
�0�Rˏ���A{��P�ky�ރ�O�?m�(�G-�P�qͮ�
R�Fd��ˢ�hS��j�B�5��
z�J,f2X�%]�t���Sg��w���T��Jɴ�gz����#�L�@�j�Q�u3�j�DY��[�{�ѓZI��L}Q�"�'M�� 1t��)J�
���09��3�U�6� 	�
�,H�p�����%�-�gQBD�azv�U�d�z��#��B��|���q��;T,#E�m���5V7ʚU����顷��8�r��8A����Ȭ����H�i}���&>I����<̌H���g�������&�3����kx/�OР�Ff�e� �N�J�(le���Y96IL��Bp�� DQ��- <��3����l�����������?�+�K._z_:�282H�%�8���0P�
\��³��+�y��A���dОA��问E��,6��oU�F6TaG�l���G]�A�Z���G�e��]�*����%4]��z��X�M��{�m ;i�(ك��s>�����k?��l���'�+�)�#=8%r��������3E��'���#��#^k��|g-��S�ʳ��2āu= !Px��!��5&����S��W����8`�h�	�XZb�~X�x�h��cz�w_O�>�����u-S˕��Ux���4���f%=<�S���j�����kV(�{mRwl!���x͋�ഐ�h��C/p�)rj���V��Ɖ�Ē.(GN��1�A���j�;&��*����5��I��b��r�t�� p�vF&a�mp s |�to&�{�5F�4>����8��XB0���W�6%�dVZ� 4��p<�Q�k¢ߏ��l����4ȥp$�4���P���(*��������;�(�Q� #z�!Ơ
7?7�kiM��>Jo�!/T�^�x�v���{�E������+�F�uq�	�x���e�T�-���y�<*���t�2ф@a����b����&�ݽ
�{D����n���
*�+�L�Q}{ߋ���e[��Vҝ�y��C0�U�\��E�g, O������㯨��s,h�I o�xM*k��JV�md4�٥7YteK�k[�!!	�R���VqP��grLfg����]4a{��7����˭p�_Xg��[� j���2C���A�zd�u!�?8�|�s7�i�_k�����HW�23.+����v�@�&��~m\i�����9%��˹j��,R� h��vu�g�����j����5���M�	�N� d����*�2~/�����U���>����?���M��hW�����cWjl��5����B��Ax|������_Jbg�cIxC�9AFDN�K�l��5�Uā��� �V�(���l��l��ꍛR�T�Ǐ�2���V� {��=����_��K�2?;e�/��7���`���ڻ:���[_���	�>�en�P�MZU�y�P���u�>�����:�9�S�*r��^i�[ gw���Ƥѥ�<��C5)�Ʀ,.n�@n@�o���g�G����,�HL��lPQBEe���S-��[9��*��}p?��k�h����l�b�W����	k�%�HZH<�I�M5	�^9��VE �H�
��D��7��ZB��V��χ<!�?+�n\g�ksmE�iV6V�eK��\�����^]��IWW^z�:ɓ�*(���!�H+�7��Y[]��,� �^�����Ot����r���,}�C�$��F�g�G��Up=�Yi�C���]�ljPD���b�Z�$r[���.�v�U}~�Z��zr*�=MeYڴ�[���YĮ<�}g_��5qm��͊���S��ZT�0	X��d���*m��D��c���L=��T��z�pc�;��@�e\]F�Br�N��	��Цh�Z���܁�*��"+m�BR�S�8���%\���W���6�C�(�"�x�m��������*l�V�59~X��0ۃ��gXY��K��=gkoҨ���$�E��pUR=�a�n���_��,Ʋ�8�s�ݗ̛{fe־uuW�R���l6ER�M�Y�3��6c̼�~�h`{$Ȁ)�,�(��E6{_���k_�r���s����$fl�@_"Y]�Y������"�/zmil�U�=	ɌJ-Ͻ6o��V�w��\��"�5�ہ��&�0�A��{�l!��ϸN8_�&��l>�8�fMv+����՝o݋z�
y���av)�#?�\��")ߥ.�)�a�	S�����B\���שp��cZ$�m����"!�8:JF�n�.e���Ã8��s��9�0�n0w���V`{���.tu@���b^�S߱��a����G��JƝ���Z���q�p�pd <�4���c��Ψ�L:���#�f �F����>G9�@��A��~4,- �xn�E�YZ����ؤC¿)�9=O:2 7�+�27����1^3JH���9�ZW�! �� 2�l8b@��F�v��5�)�/|���[�m%8bʒ��cC
cv��'ǆm�~���D����g������1�Z�v P�<.�)�Yp$0# l��74"���_Dp��spe�J"(���=4��R(�1&������}��xC����؝2��L�Q���Q�M��z�2X����#d5Z����CGA��nU��9L�r,�����g'ek}EA���L ͊��"�%u����h]�VJ��jJ6��0�q��t��sR�$�J�ڋu�v7t��F��s�/�
D�"�3��%�Y(���:��ِa������R��q�HR�o�Ex�n�Hh����㏝e&����3˄�rZA>�Mݺq�T���e�4F�Q�q� A�F�fg���ْ�:I;��X�A+6f��ނ�F`�v Lp���t"��e#(G���>�Z��ȯ ��;���Z�����-�[��.��fp�'.����dt���Nh@�:�EV�cV�ˁq�����>�k��]�#��^Јb\u�� e�gz�u|�H[�Z�^������f��`ǣ�UM�/�E���CԈ�(M2@�kA� �8O��q�ԂL '�}^���D�8J��rFW�:{�,�[N��ؕ��6��z3+I��2F,��JDVއ큽qU�foݸvUqyA�g��l~���Y$b�t6��7�i�7h��������Mr>�������^�X�¥Y��yfH�4�I�gGmI:UP`�����R��Կ��|�nV	��� ��bo��`���s��n@p�������~��%�?��E�F.6���x��������k�Ռ23���J,��������k�g�Գ@��M�џ+��]��f���*�Ύ~�c�<�L֦����������:�����#'d��YE�T��-��&��D�pS�V$�P\Ȧh
�ǡK"��D�#��/��i��qE|7J*(]@������No�� :'�`��:�^��"O�`�(??zBn^�C��!0�u�H�r�ϮN4����h�������ܬ�j���sef\�����9r�םW��h�����0���`�l_̝��� \Q��ǒ2�\R^y�S2??�Q�m���Bw�����p�΀z97C"����dI�)[=����{�&r�!�h'���m���F�Zu-�M{n1�;���t)Y��E8�����+tAD�ٮH��KIA��	�a��G#��ԡ���P�H�.��qb x7yL/�gW�Ӹ1�F]����G&���՛��=!�M�X�K��DZL��'�S�u�K
����yE5}�
H"}�@�4F,�`���BvZj�Ԉ���9s��ry��h�dVv�rX��@��!��ϼ�	�B x���]k;h���~\�D�i= �:Gq�� lT��·�@�ac?Kg���0��#�`Z=����<��9YY�O��Fu� ���NO~�k_Up�.�/_�kW���k��9{+R�W��48��Ň��9{�r��Z��`S���YS�cR
t-f%
���D��]�А����E��c�����=�υ��G4�X�̋����ʳ9X�Ⱥ� �h�:(��
��xПlT�x&r�sH9������e� ��'������G2�se6a�r
�:��)�{�$� ��K���஑�����o@B��F�g�(�Vf�U�1&N��sQ�AY���9I�&yg��u�u�Ԧg���!˂��� � 4����08�,�@����[Ę0|�N�ܫ��O
@�S������C��I��T���~�Ԁ瑞�i�N�"��	p��iD�d��>	ؔ��L�(��������ܡc5r�p,�<�~�uЊ��	�n�Yˏ�C��IP��Q��T��j���͈L;�cN#L�p���G������6
��`�\21>&@�5���� uu�k��} d�c�%��w�wi�P�0��W��:��ZA�X�QO_#����O���Ѝ ��Q�/Q����s���gedlV�ۨ�<#��e�3~{�8���WMFK�c3[zK�s��9�7k�b�]�R��S3t$\؛��N	Uҝ�m�t��8�_��JAQm7�����,
"7���z(������,��x@�23�%x�L1�44�ndO��"�Ԩ���[���s@IF�)��u��jX<)��h�-����i�&���8T/?[�ܤ�\�/&�FV?0�x`$�6r��駟�+�?�-�4	�`!-�
\:$�ٰBO�_e٨1iU+� @�=�0GA�/�{󢢨���ϖ�� �F���8/��f�[ل�z?&�"2	�CR�UhX��C����A��ɪA�3��dGd�����:	d��0�ar���֘F4~��#��h� s�V{N�VP�թK���OÔ�~�;���2;?#e�Q��
$�r�bu$H��s�K�<%���qCT*�#���[�� %'��=�^)���BVC��-��)��.+;+ܯ0Hާk3���/���<��y*T���s�pyMvo޷�:�#�t<��p\�~`�'ϥ���p퍡�֦�g"=�Tw�QO���s�GP"N�)�:L����k�eg}MaZ�f��z���y�0�,���ڦ����+�|�%��U�t�(������c!閁E�g���@�.O8h3h�&2v)���|��������� QDD����o�J������&()N!U�rQ�XA��V���R�M���KC�c��jG��y�C
F��i3�;;[�2U̲�&ۀ�|~�ٷ�J�ӸG��Ea�f�۔��g�2��5��L�F�/��=�
�������n�?fBt�,--q�VW֥� ��٧/�m��H��oL����`���~�siu��FC4�]*��./��[7YJ�>��/i�Z��F	�S�u��G�с��uAZ�zee�#)�~��H��"Ks��sr��1�}p	�M� �f	'���P�4@9$���t��j��M
%����Z�z~8`������ZE�mc�;��� ��@�	����6���U`�nh�3�$!~�`��\�f��o����Q�0�s-�I�G��)}��|��?"�D?M��\��^��h�ȌyMм�Pڣ�_�
�G�~��G����Q�6JV��7$( �fP��0B�lAJ@����#c���������4�]x5������5�̏JR�f���$_��j]7H�M����
z�D�9�ɸL�G��������f?��=N^&�ͥ�}�o���%*ۆ�x�.>�`dD ��a��GN_#�&�t��:�5��@�HA� �*��4�K>���`t1�Ȼ�NJ����C&���w_���a�q�:G�OM��J�	���gxk�~4ǿ;���aI����o1�v�?���,z= G`��{x�dS�0E���6�y��;�;�>DcPU�:�R� =?C�[���!�J��tle�2�d�r��I�����tv��i�h��Ǟ� ���C�fwgM#�H�|�N3P���|T� 8'�g�Ϩ-��G{2��0ȼ 
��O�H�KK#c��Z�ՙ�&���}]�N�)�9}!`¼$8dDmX�Q�iA�lǆ?B�
Q8h����yP �d`@4U#uh�((���c�_��: �ԉ��������֛21s� ����9�`$"�+�Um2��Ʒ�H����)8�C������L$H��w&p�@���~�R0R��2Z�3�V���䋟೿r�C�ǏʉcG8|qi�	�G�� � ag�wi|��(������Y��,�/_��G��ࠔ@�ih{�^I���zAg���Τ�ED�t�ťǸ�zۗ��qv5N�9)X4/N!x�6�/��
�ڪh�ai%�qu֨�����C�6>>!{����նln������dz�������7��`D @C[7@�/@-�0#�{����� �����ܺyO~�~[f���z:�9tu��yuVP���"/�aF'�mH���k7n�?���<s�<��SlG���e�i�`;Q���a�>3;y��|� �gL�Ư������_�~��H\��X�T�ƧS��r�=�aG��JKV�ҭ�HK��ѱi��J����	��PF�v!s��ڭ���5���P*$H�o(�F��|�Վ�7��X���o�h�����V!C��B9;H�(���s�	�Ip�@��9� &�
��)`/����d��	�2h��N�~� �[$7����_m�̵v�}0����)"?k���EM����̓�J�~�Į�Z��7p�``�Tpo:̈́��)5�
ZF��:��z���9Q5�E����Ё��Fi���1䬴nH��Ȟ��,��`$Tk3�G��u
(^��?�6:`L�ʥ�"cr���x\Wt�9��AĬo�nٔ���MnB� և���tô��3���*���=t;�S�@�V�G��/�Z��19 ��.���!P�-����@��.E��z�cc�F�JE�������(:��9�-��#�@-޳i��b<Bh����%S^�l�(�<��!�&����4��l6Og2��!�Mg�b~fJ׈F	UN��T����1�t媂�:��AԤC">mm���h�i��L-C�#��(�E`��4Q㑡,5ہQ�Ե�p�0 w	��yP���!� ���Y]����\"-ET�V������q��t�ZjX�
�l�L���I��z=LTN��2�c� }�����=f
GF����^Jeebv�亮O���F�F0��o+W��K~t�Z��кB<?�A�;���0�w�1	݌���N7��� nt��z��'y�a�Ȁ�����H�]c�<j�+�mF�Ͻ���wv���A�y�#9�����R X�<�+��I׳�2*4V&�A�{���[�w[�x��e����l��/�݊�$Qd�� yf�� �'��68ѐ���A�z���)"�n0jhS��V�p�P���x��|�������̪���k.�Ҁ:9�.�1�#��#��.Wdz~N~�WM�տ���7�_���ps�9d��"�-��H�@-�����-G���|^~�w~G�ճ���"[������4   ��cmT�2�6��Q<bm}?HP4���׾*���$w~���-�O4<�#9��&#hOn����t� D`{0K��w���_�w�=�m���7��7�d啒^;8�d���C ���݃��ܹ1=��%���/���~/�]�e��3(��h�V��:��c�v��V4 7�Ą�\yZmG��CY�C�?�����ڕV�$H���"����ޭ;��8�w�MN�P��A�����g(�zuX6J�|�g�,nn.S��k�
��IX6%�!7F��a�O�?���n?�v{%\�y(����Y���d�	� 兺��A��ڃ�D�)��ϗ��D�-FR*#�O�R kS�g8�JH�e�g
���3���+q��'QXg'Q�ߟa�2�p|�04!�޵l����7����3~�Oň}��!PR���ަ�B+0����Nhd��k]^Z�N�$^���w(Y�f�L���M�~���uQvK���9�;0;�)��o�Y@D�L2}���?�uQ��Dw�u���+��1+`�N�Ç��:�ƚ���`@kE���B��u \o��ň�pH�Μ��_zQ�F��C��"b��y���ٍ��]�V	 ��h�W�lѮ�g�0�m�t'O��ϝ��%$�}��'"�t!&Fr���.���P��t-��L�˞g"e��oJ�D� �!��݉z������oi��-:�6  {±�Ȱ���&���"d0�P.��y����h��������
Y�1���-f�B�b'��d�(]��J�g�WT$�9I�Dc�<q��H�1���G.�}��O�<k���)����^A�ʖ�����M�UPw`D�͎%2��cj@�>��1�g/��O>E��u�N�$�2+��!AxU��"J_������oj�IsJ�f�ΰ�������a;��OdL��fHB��;lƜ@�٢�%h_�yx��h�n�� ��΋	�f�@�����w?���;T�Lf�;�A::���Ai%?�����U��~����䞞�?�7����h����4M@�F�7:G��"�:,h��n@�b<R�T�'.<-��(�.]" ��Av¤�1��Ǎ_7����� 61��٬JUm��7~]���F���o��B$����&�H���R>�U��֚�Z�3u|���������8�{�����mH�g��R�eر�q=;)��.�t���I٩�0ohlX�����������Ԭ4�Mv�Q9$[ܘ=�UP�	�Y�Z��}6����'U�]P�5x�F���a�������H*�e�Wm�ۮ�.P�96R`�k��"M\.|^�ë�|��	To��Bޓ�߿��|饗�&�!����fg嗾�%9~�\�q[-��=S!{�בkw���t&  ������^��I�}j)w �)J=�*BC7)l����6�<�ڨ2�Qѐ'�4�����^�S��w���h�C�.Ar� H���I����br%D�u��tHEX ~�^��^�<W�H�eFB�R��4vN6��Е�@��"{HxXP���";�M�zA@�e�F��jLQ����G�pQ�]^]�"�1��/f�q-#
8`�Pj����n���6�\5��L�L:��Sf:�q�I���p�&���q���@���D����\��;0��XE6ɺ�/�?���pzX�fWzH`
3�L��:'Z���ѴM���x�z
���}��S��/~I�JH	��)�bj���WescK���l�g�}V���/����,�� 9��a\X8$�1�U����i ���)!���
)]�D�^��3��&���X/*n�Z�1e��3M]Ϝ�C����rx�U}s�I�+i]'�c��������#Ec�&]w������4��g������hk��#	5�������Y�v���A��MM͐�2��Ʉ��j�<=DL6K�sM</.y��^\�s��;�=+^Ē�9��9a*/�����q��)�-�y�ءv쯣G��S'�R-˂F�H�///L��[*����?K�
�S���˄�$rGٌ��,s� ����dE}>�bA;}F�I��%�'����d3b�٢:�6�f�
�dd@!���݄WLI�p_B�`�$�� Hd!C��F������9G�v}�t��M��i�%׮^ր�ɡ�Mu�P�V.��Yϫ�����b!<d�p�wv*R�)��u�z�Yzt_=| +K��l��W�� �ul|B0>�zL�b�@��k�y+|��wv���2��m�s��4dIӓQgϜ�Yd��$ �V�T	*)	P�ȽGYvx�xG֗��χbJ8�N�G�U�����䐾:��� �Hp����@�̀٢��MY����P)�d|r����d�Z�FG�đy�еo�X�� ����E�����M;��lї�RJ��nI�4m0{�"	�k u�ywSi��m,�n��K=�Ej7�0]m�D!�Ó/ʠ�&���P�1����ѣ���?-k+K��;�3
<��s�/�c'2䖆���h���	�M�#�Lg���i�u%�#�F�g���ܻ���]!6<@(�F�u �wH�|+~��H����gT�`���d�^��l�S�C�FU:6:Z �k2E��PB\����8Rl]CT�q��z\�K��pDN��,��N�-j=���-�;d��mX�!��e֘�B;���|�(r�j(��.sڞ�"H�ӎ�]װ۾45��$�L���'���qii��x
*�^/�Ƙ������r�@�{�*���닣8hԪj���7^b�{e}C�&Gi��5(��r��-y��/KV��^�gC {�p�Q��_?�QF��:�lJ��ַ��{
8sƲZ��������A�Pg��h鵇,� ��F	Ҹ������յ͕u���r��]�v횼��%=H��Y�=��:�=u�0<5n;m��H ��\[���v�`FpV)Bt"5?+�bΩ�K�V#�g��g�έA`�ی"RI��a�[}��GN�i`��pDI��
� <�s��?�:1��#)���z�ZM9|P�H�0�h%��u���2Ѥ_��\sP���?�AV|�ʖ�Zw]� ����L��ʑ�����2j�+���5��إ"����{��g۠dؑB.ke=3Ȝ�j4�6�3��3C���7�}��<��9-����!r��~~���`�n��������pj�׿�u��+e�PS 2��"���h?l�x�Q�A����wR�q�O�Y5��(q�T�+�?�z^<�w�ؑܗH8�^l*��3�I��qhzm�Id	�~JN�8*�N�ɉQv�1B ��n^ ?H<�#����ŕU��`����N�G�������ԙ� DQ��ff��~!�
=���R!���V|�(��@�ی>�9��L�[W���ư�2�������!�0ϖ~��#��\���x�牣Gd~zR��^h�m��^nW81h2����z\<|$��>�ɱqvڕk5�C���TbdR���+�A�ӨH��Ci`SR�q��q92=!?z�=�4w%�w5 �ʣ���9Ǚ ����\���q�o��M�eg������������\�zM�7t-��./K*lH1ٗ �d����}]��Q9��a益Cw8���m��}�\ؕ���k���4��#�;43���<��9y��Q�paB�<wR�R��ѐ�7�H��1E���ײ���&t%}�^E���DB?/L�A�pJѦk� �m��F���dK#���`e�f	�ӻ���i�J�#�y~(�F�{���P≩1�St�杚�ej���]��O�A6�	=4(�KS{N���4�I   Md��}8� �Q�4aY���GW���Y��Z�ON�!_`���چ���Т�6z�q� J��lDy@��t5u�[c�p_�mzJ��>;`�\^}�N�U�c�8o��u���>O %1!0�C��a:>~ř�� ���� G�s����k?|M�y�j��C���~�x�t<J~��lWG;���/g�{m�Ɍl��?~�NtzjL�4�[Z~H�O�8��k-5���ߔG�� ��/�N�(�&`x���r���q�&��Ha�5��<t*�!���v����K�5��Q�	�_���j �VSc���`A��K� ����Cj�J#�Ѝ�m��B����uO8k_3���XȆ �A!�"z�JM�i���L��0����0�Ci!=?8s�<S+�j���,mVd^#���2�Y��I�t��w������-�s�A�����˫q���s���7t��h�=g�N�8v�Q;J�;[����
�H�87�� �tB!��kk��#�s�s� )�W���>B�@�}=�/<��|������R4U�/�Rft ����'ry�F��W,��!�������+919S�6x?&q��s�aw�����kEv�$n@&Ɗ275)gN���uȻ[$�"�a�E�{���{�>uL
9ݣm΍�3(` �[��E�>=��i�R`�����\_�J��l�Ɉ>˳ǎJQ��Gk[}�2>:b� ���u��(�=��R���-��;��_�ת,�-�-�m/���&E�p� I�B��k�9�н��R[A�u�*AYffFH�D^̫9s�8����;��13~��X�*�3S�vzz�+�Wdt4Cy�I���e���ɓ��V�Hk
Tz2���VY׵���� �M���XF
����i�@�N� ��e��rd2+����7�i��^��'��-^��{��=��c~Ϝ9!�d$S
�>��3�VB�vr�.�u�����SD�ɋ
XnH�U���w��G������sO^�g/��D�<zpGV���B��a8d��F /+��2L�9*����x(aCv.	C�$�ڲ�axS�S^�f;�#��S7z7�$�"�RH�%,�)��醓��&�W���6x�!��$Z� `c�;�p`p��9��/���N
5cp��~g���#)��/g�aC���b�a���R������x�c��I��sy�D��vg�㰀�M��l�A��#!ўN�ը���S;�=�-���7,�X�=�<=V���KQ�z_	I�ۛ���#�:��>h׿���9���_�P���N��0��!Xa��}����[&�QQ������®$8S��C]8���K�d�4.����� �U5$�Q���yH0��Rkʻ�.s��Ç���6gU�7Xn'�Ґ������,��s׋��(���C&�	�dd�{6J���vU#�c�����\����W��`�7�)�dkO ���?3��:h�͎<��n���3���ٴ�\��8�|ۍ�	B}ө�fB/�(k_�6���P��4A���0���{E?oW��%1���9��1f�A�0���W��P�ե02�n�[5"Vg��Z��{ũ��<�����?���ӯa� ΞxqG�˥�Y��$���P��3�hL�sˠ=U����K�����M��	�pTȦ�|�1j > �Q��9'��t�}r>�~�\�Z�
>��|ꩧ�w�" ��/�9�� ���9�Z'!����]g�p= �bm|цȰ�0K"Q��u������2��g�g2M��D�D���g�ĩU����䅋��@[4D�0�duh�Fv�ݝ2���'����ur�FGrԣ�@���O�㏝c�dڛ�>�DcX) �����҈<��@�,�NIatT�oH׷4T����s
x&�%	1Fj�T9��@�-����M����L*`���}NV�7����@i�y��e��
r^0J$�	$�.���)�A����n˙�γ��2U���R!Z�O�\�*�+���*��+H��R[�@�%�t6��yE�b[^|F�O���ƊI�#+������S�=%���w7���-�
��uO��֎k�����������ڕ3'��;�E��@�?{������?c	��,
�]������ד���o��ʒ<�{[���or�t��������'_�{����ܻu� nZ�>�Y*Aom����E]���ɐ|�h���D��FW)���|[��"���J�
�t:=,5���j�6�DQE^0�oBTDn��NQ�m���R����D�Ș3J4���@'�6��FK02� ��@f�_xG�Zo`)s8N��)�W�Tj�8%F�+����/�"��4���z�H�;$�^�px�Iσ�Ȟ{�֖C����]�#�}F����Qci��aK�#Z\|@�&�/�s���{�-�w׊(�zud��H�x�EÚt�N8���˿�/���$��{LA�����O��'���]|F�\�)���]'��O@i#V�Mp�m�Er	�-����hiU�ݟ�����{t������}{ Q%]���]���'�?���%K��I�8��T���� g\�KW��8'�
BEXD�]R���{�6Ip�;�TL��Gaw�9$2y��d~`�Oe�d�ϪA�f�R�#
��eVnhԭQc[�����V�����TF������3H������?kc�3����:ˌӦ�jY��V�N0�� xM#�Ս])���v$��#�[QJ*
<ۘ­�h�ޕ����rS��f�^Į�~�>2��@p
@0�T2�ǰ�h�����:f,�8���K����ԈB�f�`/t �$� ��eL�#i%�$E�6,S�F�)�@�P��`L����?	���O^�겜=yBj�h`$qF+{{-j�>R������LMN�����x_fc�6>bvj�V����tۤ�\
S�p?ጃ̹��Ɏ9��KM:0d�8�Q�2��T ��s<T���J�|��m���`ie2d��c/WreY܁E�eo�pS��k'�CA%H�cԊ򭔈��S'�U���¬aOm1@
@M��+"Q��g�f����/�=�"�/l�����"����������NQİ�m�K�xl�m��G3��3jO;vD�{�]�:v\ҭ>u���R4�u��9>q�"Ui����X���,��z]�����K��;��h>3;�=	~�^�\r66�^�b9��܂V�f������s:X���(�P5��{�1u����-=}�h��Ͷ`�<'��陝����uty9��L=��E���]I����O��٣��ùm��GS)�<m�K��{��Y�z�`��j�W X�G�LeS\�O>N������w�JK#ư��ֻԺ+)�9*gO�&?����G���C9y�4�@{]��rS?�.:�؊��M0~:G^J�%���؈�,*~|�
��}-����=ir�eG�Ͷ4��*W�uo8dH�1��L�����gʰ� 3���)�F?oP�Aڻg�늎���;�����(2nE�3"D{.2�$��;�"易YF������#���&��[I�Z���¶G����(�9����>|PD
HO���;��ӄ�b6��tO��h�D�{*�T�V�ט-I�##�L�q�$����L��(Wh�=Q��
��ꪤ�� 2����ں��?�S�y����o��dF
lW�N���d<�>.�p�2�vI��ַ�#������L��$N��
��nndL�?��'����鹌�����r\	|\��-���������{�~Me������7���V�<&�I���o�3߫4�U)뵃ѥ�{��/Ƙy
22=�j�����}Ƀ$���QP����zO�FWZ�~����oC�`�5�z�wk�����ِ�wFwHKu��j�w
Nڦ�[Uì@s�� _?;�����@`ej�����ؼ�@�� 	��d��3��5NF������FEA4�?�aȠ�:A�L�1L&���	7��D]=�]��T])�wܣ�d<�I�̲�!�P���gv�\�� �Ϣ�¨�w17��?�(ta�������������)��Cw��$���X7�Iw��v��l+�*�9� ��ȢLN��s��`(��`�K&ӣ���@!+��,��4UF}�����+��g:5���a9�%�A���~�����ȵE[���)��d� ��0`ӳ1�0/��:?��E�H��Gu������I��v�m��"�P�禩A"Tk�'�dy�c�~\����-��+��뗯qXq�Ē�H>���i@�m��������G�����������H!K|
�c��7������L��c�W0y������6첻0�N����It:C�)tf���AJTE�V��[X������z-��֢������O\`�ׁu/�<T�l5du�kÒ��?p{�H�)t=����'�*�;s�<;q?A�Ƣ`/�o�%����=����[�e���W^�'���`kW��7�ݐ�
ejf^���/��ܴ������ڠŕ5;����U9|촂 ����W���Ӡ��$9 3q�*�M��Z�{
��˒ս�z�G�~��H��i����6YLo,%�"��InJ�
M�Ug<�1YճN��&z�тڷ)�@t�Xɱ��[n��f�c{��0�-�vj�)0�����8�p�%p?��O��2� ��*��b��esaLP�F���ՠO=JZ� �:9�΢:	Ξѝ2��T(�!�
��U�ߛ� �*�N
m�U�~��YH�Ŧ���*ļ 8sfMP:�f��4h��F����it���O�V&��w���{p���^}E&g�5R���]A1؃�H����ݪ:���%��?�cy�7�}HA;�j���ɬ�KW�,;L��T>x$��{T�q��076y&Ռ�Ĝ��)0����'��k@^��~u�Z����x1���@�%���̫�;u�K�Η�ߓ'N0J��U�E���QG���>�BRU������$�&zI�{�`ڧ�q��GS�U4}�dA��mI]#@ԇW��2{T�Ji��6w�3x�5�U�
x*={�,-nȶⅶ~���2ӳ]i��F�
d:�س� :��nn�H	R������Ԑ�r^
���/|���`�e� }t["`̕�+��i����@R)d0�Ip�}=���03���)�s2��q@ض�&1��"s�Z�<-�<��G��)�����Z��Ln2��Q����K�I�>��z�Ѕc�ʉ��:*p��e��� �A(@�C6�g��θF�q׬�z�:"��&��C��HL��Mb���/%�X�M���p3�ѐ�<���Y.�gdu�L��j�����!�}	�%�>�^o����?���	>C�	�#6(�6�o�}��Ayey�k٬U�P�}�n2�r��M9��L�Xu�9]O�����^� YG�H.ez"4b�o(�v�1onn���n$���
�3� Xb�flΙ�O�f)d��E�P��^ByA-�#��kx?(�BO�\I��V�4g4x�U��@�#f+{R����^��'2LΩ������n�ߋA?�4?"���>�p���g�Nhb55������1�	1H�أ�T�2��%�����*D� m�е�iP�/N��{�_�j���ޕ�����.y:�)�<��s��^�~���K��'I�A~T��L�_K�g֙�"�y��O��0�zqv��u�@N�7�Kiꐌ�&��`��a{��b�G"*�	�q�FFi\�� 4J�N��K:%L]�&2i��c��聼��PHc�؊��8�10�q�u��}S��>���09���wFT�H�fnH=7�7b��gL��`�I�;�u����iu�h;����T['�ύ�]"�J��n���u*��MƤq.�m�w�D�.]���G�k��as&��]YzĮ������(���o��/�ȡ��<ψ��$�q��;������`ܾ}W~��k����(�Qį� c�2U*a���|��O�}r��<XT�T�6E� >�I>? Ӿ��?ň1���� HL�9S�Y�@@v�yF���+L9Հ��Cy��,�N^��_��>�"�G������+TpŜ�1H0P51����|&A���ۖU�X�t� ��I0h[�M�u���5��fi�0�.�RR]ߓ�F,��z䅤�S�g�\>��p�C���mv�-�
Rz���P�a��(dtP��yY����Ԇ���W��j�v�%��GW������5d�-���0��W�h 1�W8;D��V�\"�Dj:�J��f]��s�����	��4���4$����fN���;�pG�8U�! ��Ѵ4^^]��:L���p-�X�$���;ae_�C�G�c�G���ΟX��3av"��u�0(<�b�k�վ��&���c���Jw�N.��cϷ�#2�h��՜I�=@���4c��p?8�\�9:�}�����9ҋ�H���}�h�t���4X�ry��������g��MvG�T�C��B������a�^,�pD= ��ڀJUvj����
3���Bm�X�rb]�ն��F6 6�`(���>��[MՕ��x���&pm ����U�+�Rc�l)���M6?�\|#�\M�dy@n��8Em���g�E �é�w�رc\�N{��$�����=���jl�����eckSϟ�C�g�Z3�T� %�6�t:���w���2K�`�s�>�y[����9ۓz�G}"$�����~G�~��~V��\�[]�~�gL@�W�q_����ſ�\d�-�����s��9��� }@C$e
����?)(�������y������9'n��ivB����H�e��SK�4�A��32��ЭwO_w�3ua@��U4*(����j@ii�� ��E�ޫ���l2h���h��n
$�)���!�7��k)��fl/� 	�a�ëP^`+����|D��_p/'?5)E5�ڛ������==4;+���m���m,˫��9={B^�MY������y9��)I�}�`�*�@v)Q��2B���q�֣�([5�)�a��v�R�$��o���p0 %�*X|��ȅ����2wh�"r�ZP�����A��]����ը���jV#�u�Z����>�"d6Rm4�J��%u��B�Ή�[�rQL���W�SL�#ÚJ�o$t]�uA�wSi���pJL��`t8h�~�7��i�\p,����Z�pB|,H���^S�Grl�N%mNTC��Ze�[2���K����f�+�jн�FzI5o�9���=�a��Z����v�Hao r�'8d:�cJ�jT�z�p �S��� �˰� �����|���l��t���Ḇo}��r��I&&�^���m�ڟ9yJJ

P����ufKQG�
�����|��VWv�8N���|~�S��'�ɇ| Ｃ�3� �x�y�s놼��$^��~�����o�ŋ�g������b�̙�g孷ޒ�׮������G{j�>���(�;%��h70[u~S���!8AkI�)m�?a�:=�0X�#� ��0ne�dhQ�Ğ�;F�;��:���t�	�`%r�,���0^ĥ[N�t�q��� C�
88/�ؽ�Ge&ŷ�wA`LL�;�wr��e�:u�*��Fx�V��䘂�^���߷IF�\G)����fdi���A6o�lfN���Ժq��H��/��?��G������3�>-rưo��zx[߿��`p��(�AGH�GP��j�V�������z֚o���ܼޟm#cjˠ�&�)�M�ý�1"&tf���J]��ۺ���{�:�L|����&pTƦJR�u����#�M�!����(����3ݫ�لn�o�w �� �+t��.e_1�,ۋ�ƶ�[;l�u�S����Q��s0ig���9��˲���C0��o�p�������)�&�B"��0�`)�{kqu]V6�	�  Q��O�NNN2�����⪕�1�%�.�;�Q��D��/T�߁Q&��'�����'�~���FKSt$Tz�. �T*GIed+N���~D}v}���9�vE�����w�cu�&B�B��h�3-�����j���!�e4�?�z(��s'dґ��$NW��]��H��x "�;\7O �OD0T D�8G���U�燘�
��w�X�C�Ro��NS�J�M}��R��W���`T�/}�4�+Wޕw֤�ʽ{w乗>Ev�ͻw���qfč`<�4!��}�&��4Ujv�F����,��C�k�hDצ��N�,���-�z��{æ�	������4>)�>�	5:�rj�M���	 �`��l�����SE�06����A�����Cr����6�B�rm�	s6��^}��[Ǚ0>7�����k�TN��5�3@�6j�պ�����	�����6��^FhmڊWl*o1#mȮ�Ln��7��0��V�7�4X�D���S�o���A�u�D�"J��Α�5=���XWD` �v�,1B�{��=uRK�{����'���;��&&5�-P�%F #��i�x���
�_g����}�s����쫆*��&��a  ��IDATx 叟�����~���cG�2��瘹B6��x�ءr�������g^���G�������Q2�v�t58�)���!��p.����{�A�\��������x�h�Zf�ة��|��{N��we$fv��b3�ع�`I�Må #��e��i���I��eQ�\2'��p�p��P(JG��>B�(� ��7xS�������.���8#�V+�lv���Օ:�P6Թ�ȉH$w��m*h��pIA·R�fX�	�Y9z������ #�4h�,^��)��.��֞|�W~�&���C�ђ7�|K�`^#�@vl,9L� s f���� �\��^}�eN�g��5�^�O����)�b���N�%�|q�]� pW�=OV�wdmc�����|"��H�|��m)���D.�a])���j��ASZ�qVw���c�x�S�(!;
Z>�|�z@^6%�nޱ�Nf(k�1RDw����٬Tֶ�ʵ2}�m|J����>�\�Wyް$���.@prj(�"���>��	��;�U�Ä�]tV4h�V�5�"�I�!�4���ۼv��pFؘ��TiƾM
�LK,��?K��ɴ9l_[AM�&��j․52H��6�Ds�Y�DD�;��}+���5b��լR�����<u\^}�U���W���&��R׳�g�b�C��2��v9(꘠���D`];H}��q�V��ȑ �zf�vȨ���~�舀ˍ���0�@C�Z�z�u�L��s<���n��k�_������벶�P~���s髟yEדB.��=�hE��64��? `8c⯥�-��v���N�@^�̋�^���$@�R� �uJ��Ӊ�⬎ < �=c� @㿡���(�nDf�.!m�I�婧����{w��t��	�� `�<��<���AB���~��zd]Z�O���5�`U��ݴo��a�9۪Y�А���h�lT"��U��Ws@8
o �ˑj�	�Ћ�tS�q�l�F�J��u��0�9���z#�?+��p�b���=�S�R�L�0����B#�n��-�Bt���Ƴdm���ֵ2�԰�)�C�\��Ͳ��H67VYR������	�Y� �����9���%8I��R� ��2�����'?�����J���ӂ�D��/���k+
Vf���������^__g$�
�R��St��#�	��7�7�s��4�W;�����LNp�[��bt�H�S,L��Ro�cK�.D��h�$Uk�?�1U����vz8}�<C�[�[
�3��&mYY�A�[W��#ۗ}f`��ۿ�8@���S��l�\F͸'�;�-̼^Z6�bh�PP3C>��F��NW�{�)?,O)Pİʛ7o���$�v[���� �����%�H]�	���%���,=Z����>#�#��
�!}7m���-��l��*���z���-�.�����7O���i�288�m����v� ޾{_V�B� @ϖ���9�oܔ��<~����y�Q&�q�U(��>ye({<x�,��?T߲WE*�@Q�
x'W�ߐ3G��� "k��Dr�������,�߻w��wv$a���x�(�7*Sr��������>#�D��s���]����"�Q�/Ag4	7&�s`-�E��t����tdw�r���#��/��dPF���y��.���+p��`�3i,ɋJ.8�+|/5|L8*�����F(����;� a��E����T�}'�� $Q����U�^_����K�Tj�U�����I9y�(_��E)�z��'ec�+o�{��� �Ƌl��dG���UBy��@�o탞#�y$�8�.B�>��o�v����ͧ�Ȓ�r�3�ǆLt_н��6c|����nD- %�دj����sJ��̸T�ר�킱�Q^��7��sg���C��}5"J���Z�j,4k�8������ ������T$�pfd\:a��h�b���@�>1{�k|��:��'N+��9Y�ܖ[��ɵ����ay��yv�x
J�Ð+hU�#�	:�L� O'�P�Wg�Ͳm���\�%�r@�3���0fP��B����eM���T`���A�p�W��e�x�S��-��	�]z�$��뱯��{kC��d����6�{�A�#��3�@�Bb��dҜ}��}y�K����΀ӧ����G�;���L�C�
"O(�x��	��4Հ�*j�����$�z�%�3�w����=*�=N��*H/M(H��U�m�c�9�X[��4#*�� �L�{?�(Z:�4|��hUA0���ޗ��PL�'�?��#����3�Df��L@耫�5v0di�=u4�aС���$�w���B��b06~� �"��6��ͩ���s~b�}�o��G�����E�~����7%�a�.RϺ7�;r���9֒�R3!F��i��̱8�b[� ���c˫�v��8+�/��6h3r����ʱ�{!���E��.���pxaκ��wQ.J�G��@�״���:Ɋ���a���N��K�9���-}��~pE��Yʫ��mel��z��*�	ݘB��#�'H����1I�z�WV%�edN�����6�0�0�第@z��&�uI�
�L	����������ju}C�u/�������i���[�FOv�u�
Rv�L��=7�PdCj�o=|D��n���Y>��7>����轡@��׶v%�6Ӣ�N���v��{��ik`R!��!�UU����Q������{c{KV��XC�����g�C^�x�d]܎nܯ��s 73����K|@ph:�N*Xy�Z�{ ��� pt4��y��R1[�ģi}���J1�{7R���OL}<�
�~�O*��y���)�H�'�5�/�����ƞ�O�ߑ9�}㲬.�כm����o��<�B!%��WG}�,��4T+R2[)����%j�%��@�!X�=S�)�3�N`�!ڤ�/�$�����,��Y'�7�E��0��
�b �2G����"l��+G ρ����4~
�؈���/<w�����a���P���7ޑ���<��s꼶�瞥���}(��1t�����ZK'�4�.:�Ҩarn�?K*2ndsT�'���1���)�.0��yK�[5a��(��f���Ҳ\�(fgCQnD޺tEmH%�D��=d�P��z�b͕P�#c]Q�-!�����Rn�S���!߀��ህ:Zu=���mc �4B�Ǣ�|�8ꈝt�P� 1l_���Y2K��FPZdք��qM �k��к0w�	*����|��	9y�KN�R�)O_�@��o[ΝB~��~M���r��erAl�`��>L����2�l�����Kv�Z���A&}ukUN=vBfkr��RW'��F7�U	B<���)L��k�(QngijbLΞ>�uAy ����=ܠe)xnz4��3��b.�s=;k��D�WQ$Q�w�|3��(6��g��1=5%��|$�=�|�KR�ݔrY��-��1+�l՘9�ڊ��WɡJ��1�]q3��_L�6ָ׏�����Zb ,��\S:�� j�� �"f̩(M����2ʨp � 5M�к~�K�Ķ��p-�8�6��S� 0�^�0A��Q��0�'H�H���h�:)1pN+A ���C�A*S` g�[k�ۗ�Ɇ�/�!����DV�I8p}^�~5,A=��B���~�i�"ub�;�߽��<�V�>�O���c�xdJ�����=:�Э;���
��#��{oo<�5���{T���T��v]0�>
tР���0�/�A�$�r�����l�q	�^ �"3�,.[��>��0���v� .�~�o�Y��+���sN�3 P�*����m&�9�ww�+������|G�54���2�{-�Q�'9�\�x �ν��.�Gj ��H�8(�7������5�M���Dy/p�,���:T4o ��mH-�.���p� ��\�,@^A��w�<��`��'x�trWyd�� ţ�D	J㤾��>@E���A�S �5Qٟ�I���O!&�,�\Z�S�9E�w�,=�-���u
�G0HKAؖs���fBImQ�J1gB`Ъ�4H���{
t��\[f�]P����q5�s�8�	o�����rJ�է��aBp膥�}�8�7$0`�׷نV�\�!�y=	rF�����'g��h���;o���
�����\YZ��JN��8N�Zd*`x�xf&���k1G�n��E�@`��"<?$p�9,��62[������M�ׁ�k`��S�|��.�K�:U�� ���Q����K�,�P��șz)O"r��a]4г@��"9N)��S�� �����<0:5��>��f�.#%�9!��=T���t�O���b��='DψX9��C�*���:�>�Ι��ƢEj��&�|6�S9��w��B��SA�@�����?��?'7��_�W�ܙ3��k?��&�Bq��N���@a��ܐ@ߞ��m#u���6�s��|��b~aFV ���>����������{�*%#���
�����bfzJ�|��
����~_-/�n9�jti�k}m�ٷ��6�O��O5����9�Z�c���بT�K�a�������r��8�6�t>�[@٢^�e@����s�=���v�̦Ś)�@�j�(L����pHV�{�@@�����_�o�x�W�~Gd��9��'>Կ�\�r��ei[�!��豄�f��EC�
v�NmK������G1�D�0��9���2��ss���xF�E��Ѭ���&[i�N�ӟ�3qC�Y�p��L��Pp*�(`���Xgi]� ���ӗ�R8ڻw*5����E �3������1�k
���t�@n� �G��5�����b�Y�����sa�\��I^�)�l_�|0ә1��ϥ#��X��X~V��lJ~�C��+:�p�+�l�X���:��1��+�଀a���kX�@ �O8�>�zO
���	B�H�,��p^ـ�' ׺>������Ai�QӾ�ǋ�z�EUAz��	4n��B�լ�5X�Z�;�
���h�YlFk�ֵG�0i���t"A3����|�ӷ��������}�*3a|X��&l+���,����	�I�H�k�W����;�t����|�����s ��oߺ/ׯԨ�b�S'evfD�r��7s[-��Bݻ0vH�j����.7N>" ���i�0a,<�"ɱ*���=�q �A�Pg�'Ǳ���d��ų9��$�fA�$��Z
}Z�f"A� s*�i��Ï1;�m�Y����ɓR*������e)i���r��l�uD�~31�s$�b- vE�'t>r$ʢo�šb�+��2��_ߞ1��������bi�O���\Aȅ�n�� �0|߁7���`�(��sbv*2�f<��' �@�@;�3L�a�1Q�W�}?��� S>{}f����JcA�Z�U� �S�R�sm�0�Fꍜ��pt�����X{(J�I�ό=�y��p62����XӨ����~���{o��FmB�z���*�Di,>'�ߞ��eX��wb�6��-�8 ��	(���M���6^��_���U�t�#��Ǐʃ{��h��ǯɇ~H��O_�szDn޾��������ĐO�գÄR2������C�������溂�z��G���~��0֘|��B-�ظyY�:;���-'^��1첨�񳏛�v	S~��c�EQ/'� �R�ǁ�F�fG�w��m��?�P6�5jU�M�"�����ynyYl
����8�쟳�+�[�B��B�jf#7�ɺ#�S��Z���>D �}�q8p�����׫����*_��������0�L���p-8.@� �g:�e�\6��Mv�$�+_���>}Z�&���իý�ih��eCӮ�����Eu�)f����^�ٹ	���(U8T�n�nI>���#�g�jϑ��%�D�*W�i��|�����s9|�yX���r��2S)�]�,?����<�I��p� ����/�2ی����_����?�@�;��k4=V��iwe�9��腖�u����sϽ�v{D������[����[	Q���:��1[���y���Yc:���^xF^~��z�<\zH>h.�rR�>��СY�F��1#7������f��{�L�iY��XHQ�-�5�;�N�"?ܝ�����ZR֠Ӈ�~^��t�t� N߷l*q�),Rvs��
^l�!p��5C+Tr�{أ�	��H��� ���1�4�*"vPTpj�cgN�@bHSu�"K�9�aWە˗�ӟyU~�7�����sg�r��l�-�5�t`��q��=ےI�=HX0�D���CIR�%bvD\k۠�H����l17���nd���[{F�H��?�A�+�:����#77%"�+�z(*�G��& �6=s���z�Ћ���k����p�9;h�,藞�<	J~�Qz*;BA3Fˈ�;�v��=-��3�k��G�� �ޥ���ѣ����Ǐ@��3͛Ad���Zp�{6s`��=ǆ��K#���ǃ��::Ní��@D$�Q�D���Q )�0 �P�:�΍?�7��I쨰Gʵ�z),O ����mGh7���;�{��|��8��p2�����y׸���z��q9���Qo�;BTv�$�5�3kg{��j�ab5�Xy>��/Q�F��jK����M��ķ�fta�0��������oɇ��Po��.�tՈ�o,���Tke�v��~vW�Q�<�PL5v�?q�2�p�7�}D� �����{	B`�
|@νy�dӦ��l�P̎$��	���GnG9�O����v��pB�4³���Sg�鄳���A��o�0� Jmu.��@��7n���)�����sKXr��LH#@I��ώ��u�D�ZJ ��,+�c5��:��MD�0��g�ʌ�a�7 ��]�d6�sg�P�}�h
��q���[�������~�7%�/���:ʊ�Vo�JX/��"˼d5jp@		 �:/�+��23;+��w�_��3H����/}VUfyo��{�=~�@ �	� �ː�]�(Q�T�����"�PH�@����� r� 0�gz�δ�����>�=�s���j�p\q"�5��U�������s�=��ߣl;>��@}'�ޟ^?������<˖߀>�������8��;yLu�<��M�$˸e)�\��,�|>W4=��V��C�l�������!_��?R���z-��&Nڈ�&^'�'8�T�i`�s��o}�����9y��T x�P�	W��:�R¬>������ٻ�^�G�|B��}��ʵ�g���Ȓj�cNJ,��<� �#�b�?m>����d��ݔ����.y��q�IWG�^��9� �������RŬ8}���W��>W?��8?G!�f��{v�g>���|���c"3n������l�e��ۘ�I}��~�*�@%HAdF�`�J��RG�$ʬD�$F�t��(P�!ŵ5&iiVCע��Vm��}Z~�7?�I��o�ŘҖi����x�="���?�?&���F�YE��e�G�/Q{�s �F�P� �^���@�ǣV�8'c��D�<W�T���.K6R{�H�
#�﩯�R��:Vn�'y��È�1pnv���Kj���bhW�����|da�'gd^��v�j�D��b*�2��m�a��=���&G]5v����,ES������3`-ځ#*�QceR�k���!��/����ZЪH�Ј�w���;�PI6pJ�6l� e�P��sI�Q�j�"�%H_Sh)Vr��M�x�����?�1ion�ṭ��o���r�EOo�|�Cb���ŋr��i��죈��)��N	m�<`�:V��1�D��W�aD]7���3[��^��u���r�&�(�{�˳�>��/�s�.�~�����1��/��kٝ�j�8$Sғqmk���0�B����;�,-��8-MMJCk�Fa}La�O��K/}���_�s�r��:7�Pwn�dg&�޹u]Fܥ��X�Y5�EL{.�JJ(O�{OL<P�n]U � �����~��RZ(S
<K�ja�*�(����3�;0;�Ȏ&�**^�wiL��h%��cs����� ��H������ �D����[�n�)u�o��ɩTD�=�9q1u ;�<dsV��Ȋ13"u�m���L���i�Z��h�U�9�Y-��d�x�eИS���q���Rކ�Q�
]>�%�`�'����wp����~-�������r
@֢9��&���1�������P^}�-��}N��Z��I	�lP��2$+랅��"�������4�^��(_026*�>�={�2��65����d6ڤ{'�A_; 4�yF��Y=(��3u��i�&��z������Y��8D���ƨD׬i���P;ʀ@�����tPp4&G�8��Q�.�/pW� ��1�נ�s��9�x/p��}��r��}7���ܑ�{���΀�����%�^���ī��l��bNm�%�}8[�a� C���{������{6�Ov��#;�z��ޔ'yB�@�o��A�-!I�k�/������*�i�5��Y_Z�ʓ�^g�-ਚ�ځ�@¦�ר�9?j5�(�� _�����Y��1�+�m7`zb��Ț䋫��`���(��ZA���'�mYE�K2?=)?��w�&�I�v�҈�ϩ��_d��)�����%�gi�*����'�o�I|aZڻ��{�tB���Y#�AZJ@M���#�C�'Z㇌!	\�ĭ{T\�n��Y�
����a}Vg&��ӄ̹��R"@20�h���U�ۓ�E:t��--��%mͭ��魯�ym�,IB�����Tks�Pݤv[%-�1����% `��0��"y�`�j���_��5ȴt�'>�ٷo�����r^�?�� ji��܇?"۶�KW�PsÓ"�^�[�1ֻv����P���F����}����~5b&�f�:�d�����#�sB�m�M�J7b�Fr*�_���Y��@[���������Vخ�2'�+VjR�;(	�����E���/P��6���AbX�6��VFT��eX���l�2!~���扈���.u�˺�a '���9`�2���I|b\J(U�-+c�mc���{�O�q���vQot�)��ʉ'Hڅ���� ��6X3�}�܍�ާ��[�s2��tY=��@�<��!�e>�`��� ��F	�bAr5�D!s^.YL�Y�
uF��1�c����a�v�D�YG��#zM%��� �6"�W^E&��>=@�v��|�L�9-..q� V&��^�z���̈�f�͉2�
V��YDω ?bٵ��q↜���P�H6Jv��(;V��c>������x�_��3+OQ�7c8�Y|��u�_z�%9{��3�]	k��%��
�`�ʲ��5���a�Ͱ�n��P���/q�O�`/ *�,�����Ȅ>�%��Y=o���%@Y����臯�k��b ��L9y ��ђ��߲Z5ݛB�{�p~2[8O�����f'�rS�g�~%Wus�c ��,2j/���أ��E���0�{t����?���+w󙫝Z]Z��������ә�R��`������� ���I�*7�o�!�0!t��E�������'�x�g��O����T�>p��tKҡ@�ӿ����e����Q�h91�|�K_b����Y9zl?�����4Y̰��؋�P3�*(� Ϛk��M���+]+��Ԧ�^�Q���g�*ǻ F�=	���L�*�x�.Γ 9�~��7Kg;�Aބ�ĕ��J��F@�e+�-��ҩ�ua2�.JJ7�R5�ȯ��G$���1��S7���	���A�	jN�gg��4\ȑ���$��^sʑp4�� (,�D<K������ *�գ^��`+l�f�@����Wu���'��%YՈ��@�'��3֤��[N>�tu�����@��"�Us�c��e�u���Y� qԆ�չ5��v��q&�c�1��m�Т��.� t@vE��ڭ�wS3dY��z.gZz�0��bhOA-j�v��	�9.���!JM��]�* ��U=qR��V�ϝ;+�nܠA�:&J�����=�	�������t�?z��K!/"��ǩ!�4"�F�� p!b����G���Vy��'eA1���"��q�]������V������C�l���d�0Y��7/�s�ٛ�~�E�x���TW�9NF�j,j��x �5�,3E����d�N���%��(�d�/��A�(�R}�o�Ic>6��{�U��P�>Dˑ��58+�����ź��M�xQ�>�)�X� &�|��qz��eY�s��¨#�p!۫-� ��g#v��%p�:�)���(�Z�b�,�t-�u�eA[?�#�=ݴ'��!cmq/(9ܽs��-� WႺ5 ��yn�%,)p]έR���dL9�i�M�)dK�x�ԍ|=��дJ E�W�(����K��%�pϩt}f2�Ȥ�|Kx���$8�Y/k$�L���I�Q#���L$
��
2�3��pU<C���0�ҋ�ac��#�<��0��d�8�0_�.�(s�
��k�[�Y�NX��CKs����k��:7C�	��� -ɬ\G�0�F�-e� 	�l;�bQ�$?
���ۈ��n�ܷl$xhC�< ����%����#+k�F�mj�r?Vj�����!P������Ԥ�t�~�D� 8vl�PJ���L#	� 2W��5���?��;55CP�RbKk���Hzr��9y��<��If+�59w����-Q�"��v��M���%�wp�G�ʖ�ٿg���e9u�u��i�Jt
�E7�5B�r���.H
�	�0FP-~�w���|}�@��J��ίpѐ�Ot����zs:�	�%ٻmXz��/�������z��Q������n�6��)z��njLpD9����P}��?$���r��=P��L��R�� ���b|w��f���=�.I��^K��Q��7q�B�O+��;�������RG��I��x�V7��c�Y�������g�uF���Ɂ�Gef~A�|�\�q[�轡�5jӣ	����wb6��G�n:%�h(��d`a�!WÎ�2����8*�vl����ј��	ѣx�����]=�}�vy��Y���Jwg#RCҔ=�)oJ=!���rI͙�Jv0�z �ԩ�\C��[o�� N�
Jw��aj�5f;�r��)���� �����p�@3j0M��p�����3RC6��j�g�����M��[���^f�-E��J�l슄��Z�%d�a���i]#��t�*u�����}_З�PC
}�a�d�۫Ʋ��]&����V'Ϻ�fn���Khg�Z�lIR�&�`�lS�qZ�.�^+�F��#.���A_
�.������m���؈� ���h����$~g�G����U]�R����Yu#4"��sE�q��0���Ft�!�,C�a3Jq5nlʩ�4XA�;a��>(��@�r�ߛ��ؠP�@g%��	E�\Q�z ���`@c���N�������C��un��c���g�?+��.��P�q*�_)N�a_(�F�5Q�o� !j�^
\4KEgxр�\D� �����ȇ>��q��I��Q0+�37��$�g;K3C�F���e��s�ʥK�$��,O<�8���`Q��L�,�%�!˅R��
\33�fY՟��o�%�O�3$颌�1�8��ͨ��Z�V�'�C5\$ݷ�UaL ��?��WI ?x���ʯ|�Yx���}�>t�`O[�N��k����sq��-��W������o��l۶��|�`��ȳ�>�;ڦc1k��O	f�
z��X]^a	zY��w��ߕ!}/Z�of�~3�I0H�^Rz� ��z� S +���5y��S��H��Ʋ����q��ߺ}'� ��R^f�/��}��[o�v�ٵ[
�
K�]]�ҒM��	y��W���}j7��5��U[4�0ЌX~-�;���������ɨ(��V�փ "I�$�#�{�6����Nŋ���Avj�{��w��4�l� mYuHkj�� �<@�W���-��FH7���$��Қ���,E�z��M�����ܖ�%v�p !��)HZ�L��u�o� 4��F"�(6������P�"�������2'����BDl_U���4��C�'������w�|�W>� .m]��m�>���kdl��R���A�P?X�h��7&�����1�/��#������'&t���q�ƚ�R$P�u��ke�b��Ӕn��n��>UJ�]���.+��>$��s ���K��q�SI���	�8}�T��P�� ��鸨i���+p�欚�jp�(Y3����L�� �ަ:{��eҩF�B��1n�0|"�P;GJ.0R�7^�3� �������9Ky���9Jĉ�Y���+r��;r��Y[Y�T&�I�?z�u��a41%zbv�|/,Z��kn�8R�a�I݁���M]iQ7z�>(}2*�V���fK.-��e�r1G5X���zc�g�/�e@T���"g��=�<(���)a���q�`aO��$Q�C#Mh'����@gU����;dZ��@8uBPJ�@H�37W�f� ��c���E
m99t�x�,3 �1���"z����_�1����|�u�l�MQ��	�5��B=&$V9�m�IX�q���~�!�J �O�K���[���k`�3\般���7�l��(���B6��+HkG��t/8zL~����71:F`�[XПO�߆ nvj�N`�Ƚ;Kt�K+��e������r����پs˖ %8��G���8&�BI�!23�	� �g�)���cp>48l3��^�-n��__Y��^s ��to�pU�T\�*E~���������:�����շ�d�����g(�E>fש6��N�:j<�EC�c{�q��?��T��� �+��i�8�lK6c6޷��ɘ�w�u�<گar��m�r��	����x�9�_��W�́?���)�		�Q�9@¾.h�i2R2����{�3�8��~�ÿ�3�&��S25����+�?�!9w�-��?�K���?AA:LE�T<Y[/�ڥh�
`mt�iF��a�¦��ei / �@1�A;,A���*�b���!8Z�b5�5
~m39�g�>X�J2 V�XP�1��!�N�(��_���ID*��8ʡ,��˕w����X��"���vGU#��Fh�K�ܰS��2-��cK�ҠK�\���="wF�|�]�F〉N6�S7Q�T����9=|ŵ%	r�Ɩ�\hm0@A@���z�,^�	�̈癣�,�g��~��)��_�f���c=Ҍ*ɶ�k��3261C��4���p�4��0��������_�ޒa�����P�!�Y\Kt�>|������\��<S��5�U
$\��Hwg;�AYu�0y����H9s�|F#���~iü ���o����z�d�HN�nȒ�E���(X��coȨ46n���#�@5�g_x���r����{��Miu��Ȍ\Wc��s�1����H{�3�Wc�W��	�ɸj0
.J!�����0)�3*��Z̢̦�;��Y�ha��j���q7��se��q7��Zϯ�����B�ptjB�	�����������L��)�b�2KE#�F�	�߮�5H��8��-��Y#���!q�7�k!�{#�~e�H}�Yv�7A"v�ዊ����	b6��EX���6ܬ��\�8�gB�h��X��	sE)^X#����1-���:�^jʮcje��5��UX�:*w�2�R��܌$0����7��!�W#P��!����k��Пo=� pm ��,@�q�*��H��z�����&��(W�_�)Ș s���쀑�(g^��#���(Sj���h����?���/��Z�WP
Icmv!�� ��<�a8S�x�%4�Q~������o��<x8"�����(������7�L��Vj��P~ #�3#��v�����b�|�K,/��Gƅ�(fT���
3	 >�c�/�(�v[�?�nݱS~���K��'?./����W����-��t4�Aieǎm�͵��Ķxpoر��g�����ι��/Ȩ��/���ƭ;���X����oџ�9]#d}��PE`Uv-�w����?����׾&/����jt��'�Z���-�-�&���!XZ.ʊ��(�2r��-�_�9D4k�=���oI{�	9��	޺K��,!*�5xoh�,<z�h�����&���FG�d��n��������D��$C��  "1am�.06�f����1��s�>p�J,G�}�Bo�S�+��\�`@CsA�4<n߽#s�FG@˙l�u?���a���Ј���C��A��Ӆ�]��$��"O?~Lf�$��BN���LUU]>x<6����ѣV��BG%� EӴ�t�F厚k@f	��\�1��f �����(�&7""tD �D�H$���Ȕ��E��ˌv��q�"Q�p> I��R�������Q7K��6�����|C�l��������p0RY[aĉc��W>�˼�5q .84������_$Y����:�t&F�8`n̍7�����>��%у��#!�S�L'AҲ�����=2���������-	=�I�2 ֮\�n���6�FF:gi��P��
�0��؉�Ҙi��	y�(�WԘ�0��V
+��vh�L)xD�0�/\G��h�q��EC������	G3Dl  @�ʢ�8�~%+d�P�@d�9CX�&=&�g
�Q5[�H�:����m����1�"]F�J��8X�={Y�����8	�x{����n�%��)ա.H��![�����n} �>�}/���|W>��@�͈��6�{#��m|y1N:�	�y�W0��=��$�Xʲ%������p�J[w�|���!Hy���eI#P���>d.��g��V8Y7�m�;�����xn�9��ʓlʬ�a��A�Io�6��F�Y���.�@��}��>N���'Ї�[�Ƚ�������=�w����}Eug�Y��@_wf<P�0[�����qi���,�_��rp���ܺv��+d�6�yES �a�i�ɵS<�!I'�3VPp~���r��r��	�q�*�#�Yd�Z5���Yvl�*��m������Y�3��S���6�E� o�qJ�x�I9{�<K��VY\��g��Q�l떓G3�7>>ʲO8J��#�
h�����2�;�#���"H 祔���"3�t���Fvc	p.�a�=�����	��ёr���fPE�8��~��$y"�i��"a6�$�@A�S�܊��$��o]�&�>�8'֣1����795��G�k�J[o�T߾�@�\�Fe��fQ'g�e|z��-�֦�&���w�K��i/`�P�ϕ}6V45�-ט݅v>DషYE@�kH9���V��.�G��*�JA-�����(is:����3��jԺ#�V�bd>�?�y�Ú�޽˚<5Rno��&Eo��9�I
k,���E��ў�C���̲E,�i�aͯUX'o�s}��sn<j�VLI����/��os��nωymh�D7��ȅ��v�~j�P��s%��Y�jG�����aS�MN|E���:���Vٵk�-R�����x���Q��X1i� ����8�����a5�L��]YH͢]�`�m[��S#�.ĵL��Q�Ч�툚z�ٳgi��h/_����x�a�|��D� o0� /�R�D,f#�[(˄Cd��bDM��C���׿���"A
j�I9��a�8b�KW.K��u�xn>M<i��D�0@�4,�9~��𐵹}�i�DLz��Hѳ��3� �>S�, �^m�<���y`�%�ѪN��yl�r�*p�A'��^�`n�U�3l�3W�2p��$�'D�	������+Sz �G9�s
���+��m~��Q�v���~^���T���8�F�\��lj��j����3��ȨPدZ�N����!�	U�9R"b�w	����T����֡�]�&P���w����=<Քep5OdP����e���[w
m�+=� Dw�.@��BXD	�TC3Bl�����'h�n�F�B�f����J��� �H\[�d�(�5�.,/�a>KS6+y�cc㶏 �X*H�!��!���$���m^o2U�b>O�Z�{��ɣ[Z�H�L(SLMLZk*���=A���-�����E`���e�#�G���%#�]r_m����{��{�C��9�\�uG{�t���h鐹�9�	�Yq�	�47)H�>�h�E�<� U���P/ޱm;��c,/-H�_�sM�5��]����r��y/PMO��5,�bP��m����HI�/����G������cDK_o�t)�J0�c���_�_�ڽ]}@{�<|p�e?��������M"��͟`�@#|  2� �F��o��}y���FN٘�����c�|�O�={ɭ/�k������7����B����\�������o��'�b���&����bS5�jJ��	d� �鞓h������P.�b]mq?}/��g�>�Y?��W(/������Ksù�c�Y��؇�w[k��ܩ� ���d`��_�J�6.��@CpI#$����<��ؚ:�{����|���m^��yp0�G�P�@5�$ԝ!Z��E�����#4|�@}5���8Ȍf�lD�p @�Np�p�B��bep�����F�N~C� � �M+��*�z���e{(�E�:'�1�& r,`P����
�r��5�uGI,����>��|���6=���8N2�!����K��;>���Γ +������#������j�J����	�s��in�`�����Ȯ=�	DA�ƾ��gf	iVL.bBt*F�=0^S���������k�j��1[@*��^�^x�N�֡���ԩSr��j�V�j��+}�������|��2�-�.9Gی�ݕ�@��8X�R���u�Ax�y�F�7��K͝���a��>�$\Z��7�/�Q�@MN/�	V��=��U��5���
����wc�go�����t�ੈA��s+�^��a��)'c&ZH��VW��$$&���Ǒ��r�u��z�3�s��h8��V=�M��,� �Ӳ����~�2g�9r�￢@��w�֊C�Ą
��w�C@މ^:�rB�Ƙ�4�kfXj6U��3n�'vŢ��`���;Bk��QΔe��hC��O�?
��kpa�"�A+�ԡ�#�R+ʦ���푇w�J��BGݩ `��-���H�.V
,��n�Y��%��Q���3\ʯ1��"��!-�k�޻k���S�����QfTp=��2�J��$}]�8�TnP�-��_	�hۏ����ڵc��yyq���/�5.-��};;�e�𠴶d���g�j�(?�6�����_vn�"m�F��|>L؆T*�D�WȭJ���^�|M�g�lr�H��sz�(�u��p�1f�a�V�}��2;��e�y}Vv��-'����\�uG����*�"����8��Ә�֎�����B�*�N��Ժ�ut��1󶢀e?L-G�8����c�%��{sc6��bYݤ���D���%���t=!�D#�e����D&�8y������-��:;'#A�V.����w��T�:��^^��'���6�"6� ��LV��g=KI����ߞgN�e"ThC�j�����L���F�} �L7�ڷ�>-�a:ڻ���V�M"Y�����N:	����c�L<%�}C$]�s���α<�ōa� ����IǨ�
��Z �P�4-� ��H
�N��k$@a��Q�zOg�u��laor����g_�Ғ���+W�XR�����L�aP.�D-��R��Yf��a��tb��w�v=,G��%�LA�J�A�Z��D��F?C9l7 �x<;L���c�'�G���c�+�n3�Mb]�$Ѡ�!Y$�Z�Nb�#D[��6nK
� �Z�M*ȹt�2¡CGd``@�z�dێ]�� ��}�{�>[}�RI�b���MN�[ ٶ�7op 6��k�9�E��F�c@^+�$(_]�~�u[ԁ�� ��ۺ� �#��r8+5SwmL7�
����>;<�@�t-��W�lL</F�%^>�侉������l���M�!�ar�:fdj�uS.Q�/�"���4dM�)�|�:N��J��d�s����0���q)���*V���˅�6���
lmf�*b$=L{�=-��S���zY+��ua�i�X	��vf��ӹ� ��AUi�E�єr�6�rlr�����gJ�ȸ)�O�=T�yQ�Xr��nH$	�(���}� �d�k��=���zg�d�1��fk+�n�T�	f9ޢ��z�&��Ye�@#dpUr"q+u!��L02�E)����;�d"��e�Vܠg����tv�����������PJ�RT���ݻ�����//�47����}�e��WM^�J��q@`r�(ag�R$n߾u]mu�<��I9w�2A2��T@V`=�"�C��w�J��pb]�z�ۛI>'hTpY���!:�嵂��_T+�9Ѕ����}�$��R�@�ea ,s�6 ������s���Ԝ:����	���#z&��3� R���E�UA�@{���^/���O���i��ˠr~zJ��:k �#�T�1����[Y�KD}� ��B�6Š��.BJa���Z��՜��>ј%߭��O�h,��j�w��oӱWW�s�xm2�����u��_;px�l���҉������+�f�&F���l�֝##�����J'c�h?�YDH��p� �'�Dmv�?���],=8����0�O�AA*Y|q�:B8A�������H��V�z_VQ=
�
^�X3�L�56��;/ɩs�	^4^ӟ�B�43(Nq1�Ή�Qˤ�Ȥ��Ii� ��~���^�gk�l��j���! 	S�#�ql;&���u5[�;���!=����"��C�"yq��ee='C���P���>�:7�$ �Օ^�c�Z6��#q#�x�0%mSVqM�;  ��͍k �G�?9i�W�7 �r�q/��F�Y�q'�M�f� �Q���l�>JA��g����
UEa9P)9�N��ߕ[w�Ӧ�xL 9Ho���+G����w�}N/�l:����5y����;��� ���F�����p�I��
�+ds X�}(U���5G�0��tQ�oḭ�F}�FR�t�%4h� ��$ר���@�wk{7�05!�:Q�+<;�8�Y5u�� A4�Qb}/W佯��� �`nS�A �'��s9_�l�����~�yf�,q3bl��KA	�}x�!�m�"���d=���C��ĸ�$p��),��gM�7���sq��	`�1���Z�N�����48�
�f�_Xo��k$����4j]ٖ6Y�g������&:���*d�i �I��rX�j�jc�|[d�X�CA�xԕƢ&Xf�����++���g�������,����vI�^on��~^Y_av2�h��� ��MӲ4;�l��j�L�g�0?����kl	��b�$|�fٽ{�L�NrL�~u�(?�~!��3�ξ-[d��t��(*&·��%Y�}���[����Ǉ�w�ɃC6�a)�D��YSA�������y]_[#'º=���B������^ٵs�ܺ��Y��~vR�R�s}�]$�V������� o3��	%Vhv�y�ݨ�n�V����[Im�c��٠�jd4P���4�R�GbnSSB�ˀcue^�ȶ�-�ȪD�/�ͳ�i��-��j!/�[�8V&�����Ӧ���(�ʗ4(����VjS媑zV��, F��\�4:QF���� ^0d6���t���n��Ǟ�����^<ܓ�i����]��_����ɳ���>����z!WzQ�e����������3wvW���G���3*Q*���.}/4"֖��L:D�%Ѝ)꽵bL�h��Jg锊7�F�ț"�������B~���g�z��c�U��|p��+�ei�*됊��ڢ�<V7��F��P@kpCs�<�iX3�7�V��6�(Ŋ��G	�х#ЂOQ��q*�������@a�ڲ0��Gɳ<�	sH{�(>���p��A�ǯei.�ה&({��G�ν��5y�.�=t��p��ȉ�l��l����YD��4p�Śm���^�.�>�ֵ���Kj�j P68{��_�jnm�4U2AG���3�`e�4+[6Ҭ�"D������U�9m�0C'F��,˸d�N��V1�A.�#�Q��۾��,����< �N�2>1:h�z"��H��1�а��qye#ׂ���ۣ�����|~hg~���e~qAn߾ICݟ�S7�G�m�Y�P�b�ŵ�"kC���X�@e���; }Ͽ��E��Ƕrq3rP����{{6pR�^�T5���'e���TC�2k���Ize�w���)K�g��׸?��B���oz�2�3W \+1{ aMbq#^����edB����\'�l"��s��J���܇�F&�r#�'��p�`$���%�*�4P�(C\Q�1#���=M�w Z�z�[ZZ\�'���D�1g��5B�k��?Q�	S�޻w7'�NN���c6�|C��\����^_FL��tu���&���$]��t��%�~��zYb��Z.�.H�~��(Iǩ�d����Ųl엹jA���u�0��^u��z�_?����O0o� �-����_t��,/����WJzM˳3t�,��}��Lˉ�G�ȱc��?�
[�! �qR%w
3��9�6ݕ�l�G�<#3S���8dS�3Y�<9|p/;��I�3s0�A�?�̐~��m�g�Ho�A���W*���������g9>=%= ܀{�rF����4��r���z���W�̩���-Q��Tcu�g�[g�M�W[W����;!�f_12���,�,�rSAź�801���~=#�Hnޥ��YKv	u��;h�"�Ϗ��^jN�8 ߰Z,�./��ٽk���o����g_X�_��~�s��{�A�����o�_�V�;6��R-�	j����*��%��M.�g�>x2-%���D˞Gnht�0D<S���VO��X4�vJJ�z��j�J{�Tf]|]yTX��Y�l�g��%����I���/\R�9&��3r��]�C6��j ֋֖����jQ�S���Ь��'IN���`�S�Q,(�HbTZR�-$wҰ"+Q�i,I+�D�M��Ѣ��&a��r�u���@���Ȱ ��%ĤVl>+����om�����N�0]��'�$C�Y%�(���r��yɩQ�3�ȏ+�o��u��`�e�τq��A�_�Y�r���>�����2�A��)�6�u�H�'R��Y�r�U3�Y�U�Qã E�IŮM���)�1������w�
�vb@"�VU���9D8�j�Jgy�����t�I�(Ūl>Gq#N'�������J\;:	�85)�bB�
����{�����������K,]�tQ;���i��O��d�������>���z��{d�|���&���-��:�	/84�u�.���y��P
�^�ͬ��@���z ,�H`��E�uN?����@v�f���`tnUkDG^^�o(ˢ;���]�S���b=k��� *Qп"Le3�>K2)Wz�-@֔���P#@`�kϵ{1�R�ggP�]U�(���5voY骁2a����im�A�{0��P�^(�mߺ�D[K3�)�8�Y0�P$����w��;�VQj�h"yz@���B�����l@�Q�A.�Q��/�ȳІ@��⌞�Y�<��I9v��:�t����V}V���7n��>�|�S֝��o0�������5$��������e��o�H�Č�qD���z�s��l�mC����#[�=�L���5��l�ɞ8�(J�$��3�8�WmP�?�M��1�/�N�K��y�'�mB�X����E!Ѥv9�g���M��fdk߰$���d�J��]���\Q`��X*ț�F���4 u
�z�1$�@ޚpF��F�'���mK?[�5 n�`���e���mi��+�g� �ꨚ��
��1�����!�kҺ�E:u���Q�]ۊ
���"{	Bt��X� ����-(�MMNKK*��d����V�JN�J�
�H�81Bح��Ҹ^#�"��Q3+ͩȻ;��|��ſ���,����g�z��Ap5���+ŵ����³�+[(G�l6� ��ŷ]��
�3^8P�F�6�י�Q����%���v����K~�$����Nխ� �A��M�Y��洢խRV�t��=�|��|pJ@�H��F�U������Mp�WOK�#!t�a-��� j\�*�b����H���������=�₰���l���x�x�~�}�û����i�<�IV�#~^���g�Я���tuu�1lû����7NS�F�;ݮFnA��-D�Q��m Gż�l�"LZ���ؘ��PF�ĝ09ڋ�"}Q�B���'\�=���Y��>�u��U��S�����sN�o���M��Q��۔��� �Sp,\Sȉ�B��8���6����(m����?(��upfv Z�R�X8GD��١K�69"�y�ކ3���vz����@��e�C���x}�7���׌���^�)���C��?.3���I*���r�H^�pu�9���>T9I~$�Q/Db�<�瀜(9$�"`���-�h_V@@�[�o�#�C)��_�S�I[���c�j#�b��~�� ��Y�壗���#���W �ep��hs��#sѨ�<
@���%��g�,�8>>�{�d��^9z�����,UVQ��������[����C� �/����8�� bg�9F���&R��XU���.��\^rz.�(aꙪ�cj�{���)����y���oߐܾ3%_��efbT���?��I��o|Nz�;Yg5Z?�s�ݿW��-����D��������!�������� E�A��}���%�I�[g�e��k�"PŻf3Z�5��x�;��uf���,}0�Eo= C[��3q�V9�;g����(t��,v�w�N�̞UWʯ��n��g��֦�V�iI$m&���ʌj+��>(��������uVV���X�C7�Ơ���o���y�ˋx�z���f���.ұ�y� Ev��A��]�)�N�y�W����Gu����M���^�y����p޷oߡ�#�xפ��#'�29�6��nV����%�4Ť�e+m,��C?+�����S�v(��pU�VlzJ2}�/��8�!�l���^�T st}E]}�m���_�����W�����u��*o�Y��^\�ӿ{�����G�?!K
��v��1v��͛x?����D99-��ċ�ׂ��tD(�W��:�	���R\_ �=�Ze��m�|����޺��djzRΜ9��cZR9.9h\ ����xL=cDz�u�wS(�L� �!{�Q�W5�I�ٲS�L��k%�t�9W���Sn?Z��:W#ˆ�B+	E��]�'n�}�:!���kj؞{�I��G_d�Ν��8����V�8P�/~�����y��(#U�w�l+ES�eB� bܵR�W
*b��.�3!����g���$gֈpX�O��(�=�q��I�l+�s'@��#����}`�
"7:V�x̨Ԩ,���cUs�)���=�,��Y���-ϵ�1�o m
ǜ��n�dz�h�U�ω����ϸWD-����X���)��҉f5��x��5jǜ<y� ���r���	�.� ׋�pd����8�vf��l�����O�8�)�:���R�:���VaM̸��v��G�Ro����!����� u�釰�Ѩ�x�Ȏdnݶ�5��,��π�Aw ���� 0�.>�5(�a6����{vʁ���962B8���_XZ$��;�?�$���W$����ȁXר�ȁ���:�UUo)�̯��,=~�|���膌F�㣣�ض�wJ�9+[[ID>��@�J�B�Dס9��6�t� #�˩̺�֖�V�{GK��2�(y,-γ̰S���z�X�&����[�?���c����7�|�D��/��#�ex��sZΝ;Ge^q��բܾ~�Y���^f��H!�*1�S�ߘ��HF�o��7�J�e�Ƨ�ɥ�����K���*��d*NM�D*N'^�|�u8��uH<�"XE��fq�����g,Ӫ ����
�*j�������w�\�Fd�z=jG�6vEL�xQ��qut�ʥk��b>�M��{&�vuM�?.��<������6R�D72������흽253���
v����{�w٨�ڽ��<���p&P��Ҫ���JHcS��*��&V��O����;��?��q���ש�y}?�)5����OV�#�k@�N��2�h��So��XmT}��A���рM8S�>�kˋ�>��?���=�.�H��v���rc���_��V�*���#֒���j�S-�_��F+E���k$ܡΆ���t&P�J����(���G7�>��n��
[��tc����n��uq^����|�~���"�i�0@K7}�n���>ݼ5�/�h�H��9BN�}�>��Hl�},��;��p��8�	E�j���B���$���*:�`�X�J)j�*�?��	y��'��G�#�BExt����і�5V�IF��WiL�-@	�]U����F�A�*���j�b�lb�~&ůP"�lP!�D$�3s�О�`6(�bI�x�YgZ;	.r%kTEwF�M��D��\��¤ �擯cm��tȸŒ�:��L&��}���L��v��8Jl�èр��gYY!"5����G�{��(�� #sKN����G7�|�M�N�\�@�2�G&�i�	!�������u�K�=p����͊�o8Bh��=�c~f���W8��>e#��dh1��R��2
��R?�i{4�f�9��������'���[w����R�h����a���Rf���/P"N��@tUa]A�6@�62 �s��f��;�Q��41���X�	x��s�<��cҭ�PoW'��@�G�g�!���b��p������!C�}R���՗_��_}�Y  h��x�1:���l�2�!��ؙUG�4gW� �	/}���\6%���>����cz���%��F3��̆n��xt�aZ8J�ȅb ��ĸ�t�3�x��>����y�=�_�� ~�9���;Ң�sx�^ɤc2;2+�umQ&����t�����Wp�"�x���Pe�,��<F5 �XZ��R��g�t��r���L�.��U7}F3�R,�Q����s�vٵg�\<�r�	�;�l���fy���M�����k�J?UOk�	�pkt�Yph&�w��X��b�UI?���G}G�|���)ǉ���8( ��,/:�t}kz��5��=�k�:26ɮ�R�@�W��(7�u�k�HL��2c`��m%=; 8+k ����}W��+c#d����p�^D��ǁ���w��9r�[A��\�Rs`�Ӏ������G��f	�`S y����Yf�zY]�Y�9d�rӀ��e 
���K���W�b�馔��W���8&�ȯ�==S{w�����;�5�j=U�.�X�V��A$���E*)����NkD�ֳ69����+t�M�V����s?9rGVt��h�Y<̷/^�E�s�>��ن���2��d5_�FH�uӫSh�J��6�ܥȿE���)��t�lL:��f�ʚX���P��^���i�U��-%�P`-Z'Ҳ]�޳9;0�a�/����o�@���c�{�v��\z�"Ө`��a.��Ƚ(Z;[�]�k�핻�C��gĵX�3F�*�0O"�H���&B��B���U�v��A3�ah`���q&r%CJ��6���?���DC�J(��87��4�"O�"���h�B�(f�h4����Y�d��?X%)���^RQ�F��J ~K,�g���z�N2!�G�O�M��G�#R�0�I�'ȳ������#�n�����ш���ݺ\���~}m��Ѧ94��������w�U�V!������^����W�c��n~8�i]?l#����Q:b�w� �@´U,���:A�����g����C9s���&F��,k�.�b�zr�P�	�'����^�;D� 0��4��Y���Γ>κM��'U4���^� f��s(�|751��G7K�����[��Ɗ��w��5� �3,��5��#;�n�ұw�o��5��� nq~�����ktR)�ӏ�_��Gf�1��g�1�9�ΐ���?�����g��#�HK&���&��[�,�/�j�>'��S<�X�XS���}�Vi�yl׆�G�_�^,��[o�&���G�M�d�~�}���@����ى)��8%�@��m�(�uv���ZQ��*��y��y��2�P��蕳/���>:�$��u��pF<��
``C�{�to�r��m�N�1��ڮ�E�=��nɎ��eiyM����ud��{(��y}�o��(;wn�8ۍ��-HoϠLMMS�3�A�{���kV�Z���I�x~�@w�p��./�+�=}ҥ@&���dr*lMO3PðWd�AJ��
��B�!�>u|82N�|p�N*Fߺ�P�f�(`C�#VZ�72�Yu�H߸sWV�9,���P�T��,��7e��Mvm�{ӵmΤeq%O��j���[ylU��%2=j�0�	�|���Q�uu�?5��'"���=����������N�+}�򃉛w�ί�jA6>!�F@?k���}�@%��q>9�_u�̚�&Y���9��:\��A���VgdmqV�RN�g�����%9u���������Wo���6O}}�e5����t���NY˃�"d�Cs$��+A,45�ki��q�#�7�p�ob�� 0�ù�^�L�R�T��ƢQWn	U�"���n�A6I��ր��{�!B����uit=k_���ԨmZN�q����Ԭ	A�*nz�ɻ�0����_=��m$�V�9�E}7@�'��^���3/E�rMH!`V
���̛�=�|%��u-�@$^s؊�}�ϳs
��YvcN� $�)#�Ś���29���ʈAĉz%.�L,�L-cB�ěx���g#�ӵ�����1
E")V���s^?�����SG��Z�X�����Ǌ= �Bꌳ�^��b�n�l�{-�����?%���JC?�d�cA�S�ef�©��8��*a��������
�(Y��QnC�|[[33�ϟUP0m-�S��	��\K"4�LB��ҧ�$����yu$��y<1ݳ(' #˽,&UoZ@�zI8�m��R<(�a�ܽ��0S����7d��]$e��:��Ρ}�e�:p�0ejb�IpT�I����"�+�݊��~�!*���u�����eY�2�I�Kc�^gN�M1 1��<����`O*H�l�+����/������ԯ��`7��i�P��&ȱ���5z�ʯ�گq�{�1ez8�;����t�y��9���_zJ�me+paU��ۧ	�R�Ƙs�̥����E��&Z҇z5 j��7�%���l�Gd���>-���V--b�V���M

��H=7G�ڦ�z�C�ťy~?��?=���Q�t*�X� sLmX5��mJ�42ޘ��lÔ���J�@�7��ݣY)a^�I���%�T���Z\���A�[M��H�ϗ����ILEP��@�C����"�CW�K�Z�..�$:;?�_h��k��4�����{�2䡽{%��=Aa7���H�[@p�W =������4�w�4�A+;���%�������U�dt�s��(N�y�����)�w� ��p#�QYݲρ���h��K��{�^��5�۵Ҟi�=����ZM2by~�+W���j�/P�K'�l8�����ϰ{��Q�;z5D�AhT�m��t7����y
�á^�&�I`�|yY�hL���!���L"e����Jd�{iu�xh��1i�|����r+�g��"�:0<1ycfTL~����8�(���m՘��Ө�,PKg�1�:%Dq�0�yӰ8dZ��>��q*q�|�8DFTp�-j@q���?y\j3S�p
�b�Ƅߢ<1��g}�:�x�����rb|���=�0�Arh.:v"�`c��+�r�`\?�H&<�I�V�|ٕÒ��Z��x�T�"ex���)���3o�o��
wA�{��E�Bl,��0uXf��U0�F}�5������+����F++;9v�ᤱ�MMt�j�@f�l���\��mq�J��(�P��se�A"�2��#�nzm?){�7����^���S&B� ڲTs�
����+b���<O8Fϧ5�'WJ���&i�lc����:B#"�LP��8�a\�]����q��%v��?w��ߕ�%��WWW8���Fl��qںr
�<��Ӎinn%?����Z��{���+�QIxqyYΜ;��|��	L�F�0̦�ӧ�L�ȳ��������� ���O~��%A���{��k�,O#fgg���:���}$�6���Y@�	م���\~碼��o�t�����f{*ʋ(Y�J�۷����)�c�࣡K@�N��}!rq�i9r�]����#w�&Ű�R
J �BK%"����TI�,��� x�_X������XXZ&���Zw����;�4`Z�dw<<^xo {Ik
6�O�l�Ԓ��w�����t��U<���Mٌ���dA��[�_���u^������[w���,�-����R�T#  �X���p8����G'l��� BEW'C�؁813��8fZS�k�����,O������p?��:f�A��<|����(@�}z8���2� R��q0�~փ�	�Wd3��3D� G�?�g9� T�2��Qfq&8�6�Ƭ
���ٙZnij�̔&����?֫�Ұ��N4������t�ƏF�qړuY̮n詿���D�SK�4ko5��F"��(�L�$����Of'4bZ��M��R��"���M��1��)���!���dǥ��F=�]�'Y7��jQZ��HԬ3�u�
�8<����T<���CM��)�
��{���1[q7gĢT�h���1t<��g�J�:/��>˟�1���݌��s�A�H���́	�f,�F +H)�QT
��AE8���2�8���LF@����pIi1uLd�� 
�-��,F�1F5����'�l�W��R��%�. Pb��Sz���N"~�����is�x�2]���z&tV#��� ��8h�q�A�J;v�9Rag��b��T	��i�V�jX���x#;�`�$�,y��\'�:�0N�޽2�6b�)�����Z��8�R�:Y���_�{|�wo���w�<�=?)��c�����1�	�~���8��//�N�-P3�N�1h�d��}�'M_��u��Ǥ�)�'u`R�P[��`��[����0�S��
9H�#�IN�zC���E�P�Q����Ѧ���>��-[d��-��ۿ�I� !()ݸu�\�e<,��j���C�r�j]G_����)�T j 6 �����o�y�G��G;4^ �b�2:���A�g���� w���  >��������������q	�pBS������`�BhC�$�lM�/�������i�%]�;z�{w���n��z�M�.C��N�aN�#m�����8���A ���4�AbD'�l�"�+�*hw��T K�B��k7x!K 1N��8�,�����-�|#c����횙��sxc5�>4WW%��H� )4�=N���;Ϝ��*f���o���m�b7����Q�	Z��Z��ş�b	m�y��&�p��	E�N��<��ȑ�q��E���0/�Z���a�B�J�^Xr6 Oͭ-���U��Z�w�^c�
��9�`̧����tS��C���Q�I���8�<K�`�b`}��~����~������b��y"j/�gr� �1ј8��CR9(P!��p��ꆊ%���M�F)؄$+����.R�%��"�FK��kl�?{8�iL�J�BM���K�.C��c�D�i�㟘5�������x���iBէ��	�)�+�x�D�������HJA��qs&�Y �����!zWcuYT��T�Qhӷl�%�� �C� ]r��K�CS����V�B��"�
2) -�M���j�d�HԐ6�6��L��C�F��X;�&�,s!����;��� !�;l�L{�5��*i�O�D�uO��Ci~>7sو@S�uB��ϝ ��-�Fd��Q�bt� Y~Ą���=
W�0`���0��oQ�uDz��pp�" ����-����%��r��?�0�Z8`V�s��D�N�p��δ6Ȗ}}�R���R ��n�Hn�t��"*θ�V���ϐe�|�N�9	��`�o�m�}���`���7�Z��s@�"
�@ �-�I[S�`\�8��Ky#�2�8#��>��^p.0�!Ø
d.�y�҄�2 ���"��l��t� �)<]+�?R���\��u+W|��&S�Dɨ������O�)g�:#�s3$�6j���@�&����[��͛���i=z�g��?�m���y`�'B��b����dx�����~�;�"ZSg���k�V羸�ƙ+�-��Tk�q3]\���*A3�X��۪��yG�s?r�CHSM켚C�B�
Kkr@?�ȑ#n(��9pXv�>@I��7G���)Y+��=Ю��&�\�N�m.g����%�� ��
��O��g�v��C�QE9A32I���!���yXn �m�u@�a����e�Vv��lM ��
�3ٜm���i:`��#r
V�Iɯ��@u{hpX���'�w��^}S&�gM�;%�K�
T���������oF��~�{��Q�����sϓ4���Jy\maSK3�}��
�ӳ��' :}�טjl�&�T�9)���ޡ���*�cf�FF$y�PM�{A��Ӹ�����ߤ� ܡ}�Iwo�<������g$Ӓ�	�W��Y.��uo��t��AJ�Y�?|đ�'�>�L
�FU�[�4c*옰��_	���?Uy����k6�D8;��=ZKWLg�Oz� _���z��6��t=g�8�1L)��RM�Ӧ��*5X\��Mz���Tkh���M�Ō�r1Ԧ��
�4��@�՚iz�"CAdNQ+3ܘ\��y�	��i1˴x���{�"-"��(����D�%�Љ(vرR��]&	UH�F��L$� HAYY�lD��~J�y�Q��j��;v����:vR��?$����\��)�`�cJs��6dt� �0�!TM�����lJ<�U��+ȉ	�2:~ǟ��qʰA��S)ŏr	҇���$�!�G�S�p��O8�jk�ocR��c�>��"�u� D�)�2��@�w*�#��B�6$A��E����٠#ȋ�_��+_�͉!:��.�w7B��Y]8ap}�Mk���q�`4ҬFcQ�k��)2 �bj��P���� rD�y-WԈk�Y0�Ζ!KnD�������ճ���~�Ǖ��`*� ��ߨ�\a]�]I�=�L���r����o߸M0a ?Jp�	�Q<�?���u�� �3�k�O��i~�y�܆�~<e�tGB�f��'WPc�sv��c�<*J�$���xve��)q�����M��nH�C�S��tBM�8�S�K
����������[�u=C	n�G���7��1/*�2�g~ZI�mY�ϧ�F����c���O=#{��cV?�ri�� �/�^i���Qg���⳺.B�=r
�D.�s]������{� ���L0�{�]W{7��0� R$@�A�F)Q�]R�VZj�tڋ����ؽ���q��J+�J��IQ�� 	Z���w�c�w��U�]~_���@y'D��iS����~�_f~��,^^���]�?c���"'@�-�%���H^��%*�R"��NIL��{�c]>,]�db�V��� �ڨɉ1���n�P�����X����|�Cҵ�q����W�'�C�<?�S�b(71�9��dy[7	��Z66�o�G��=����������#��- d�'8�Ѓ�;y�����"�EV{qR�"Ⱥw�y�}洼��o�`6/�>�4KZ=��hF�����~�Dwd@�!��4�-���}�9��������/Q��d���a������ޅ���B7���S�Y���\^^��������N�lq����E�Q�9j&���}�Es�>��B�*_��W���M��C/��xWjg#�N;���u��?��H��-6;�#x_n�/+��ȏݞ���~� 5� +$u-��uB�� ޓ�`6뮑0��)��{f�Q�A����sm��gnQ��J(�X��B��vj@�2��u90�(C�;-���<�!8H̆��!:~�J�|('
�Q]N���]�b�����N�վ��E�����	�.f̳ۂ��9y�gX��[�B񰝻����{�1�S7�:��?u^^�
#����r����k�L��NHˏ�ܳ�U#���Y�TBYq�����AھF�e�] 8�t̉T�-s$�¡�l��v��e��`L���������J���[m8 @� <ǃ��;��(�'���]�ԏQ�  "td:m�N��J�ߵ�1���Z�R`|DX�hZ�[W���udym�����aZ�H~T��o X�a����uF�nȥ	z�ݥ���Ϝ�_ �m�����6ψkR��Jx�8�0P5�Q''5�D�zQ{g�w*K$@r]X�}�C��A]Sz�7�c#�� @\V�n ���"�����}�k
�,�v�E�R��]�5�$^��������-%D�����s_�`�Z�8]h�Ex��+r�[�#�+W���3�s�:��{A]#}N?|�)��{�K�fg8&!s���s��67婣��^��,W����8�`����)��oj���b�G_xQ�򵿦���vJ<��eL@ן��z�db����<sV���'dB��d�+[T�>{�<3H m����]�,���_���g{��qi���QP&��(���O}J~����}�W��~k��7}��.��'�q}�@{�"j� k�i�dcP_�����G���ѵ�l�lT)��k5�M�#���"C��� ���������7~��[�φ���K�(��3�	�:0�c;�W��D6��G��<����[�z�<�����{�&Tj�ǹ�!f��Ŝ:S\G�i��s]e  e�5a���/ɭ���R��)/ ����9Z�a��E!��o ����cߖ�����2=;+;w����-5����q���t�pms�6� �P|��?���� ��0�VOb�5�j�ҡ�r����s� hU���U�TJT:�|��G;(33Jd�����:�~�`u}-HG�h:f'��=�E�u	R���w7l��j���
�%��A�|0M����!�P�G�|@P�s:,����i� �#6놜�:=� ��:LYa����(�?(�V1�qB�䏛�R4�5#h:Hfī� ���z������$焑e��)��z14�)���aI+8���b�%�/�"�Ξ�d���wA�yؘ�`�eB�&2�.,/WT��DĆ�lX�4�� Jw���tµ�,���j��i�h�+�!��ǧ�!e�>I�˒�c��~:g����	�6|��kE�%$	BQ@��5y���E��5"p�%�ِJ�Jp�����:��M��`��C�0�hZ�t�Ԛ��r�X>�����,_�(:��m๡ke���q�DG1�A{~$���BF��@��k#ޞ	y��Vf嵴U^�3,%9N����.!'!J�!�
A(�^���!�	u�q�R��ᙀ�P�3qr,+$6wIZ��Q|
����Tk
�=u>�p(�!��-��u�9%SȄ0��a��9#%�2tln��fu�{���c�z�[����C®#O�%�7>B����A���;SyW��)���Uy����
.�&'���������ۚ:u\��g��2�`���"������ڳ�[�1����<����G J��9yH#odr��ט�`����=@T��j�C	���ё�� zM�_~�+$��3�c�C	���\���z��s�y���̗B��f!���L'���j��eQ����1p�(Gc1��3�9��g�D#���q�h�xh�bT*e>�tƆA6X�W�ڔO~�<��p��N��l��`�0��v�	f([��������AQM���/�=��� ����p�f��b�c0��
���V7��V>DlX.�\�?��OpV�> �>x�Cql�[_���S�63 1�5f��~�g-��k�fXd�{m#��cc�lM��!�2�^����!�S�Ro��e؀�X�<6�:�=�M���=W�^���*�Z��l�jx�@�� A}�����V�#?6?��*~=(����j�I�I�cV�R9�E��)ekS6�Zʻ�{/:R'::�뽸Km?caC��j:��t:F MGC���Ji*b���֡䵢j�E_	�:Z����ph#�0K�8���3�Q�����9g����!'ԏ@��7��t>jӸhN�q�p�����4���F�3Ͻ(W�Vdtx���Q0�7K�'�ȇ[{)�����Q�slzQf	@Dd2��ԃ	A_84j��p,]n�k/k�YwT[�\ksI�78j�H�����b�� �ǭ��@�$�� ��_�9aU��1�䡠�;r�#$�(�nM��VR�-�F�[�6	�"� F"7Ʃ��F��cɫ��9b���3a�<XG�9wD�L,��v�h�%+)z�Q �gNF�T��e?B�D̀v���'ym/�2�v�� Ԑ�eƔY>Li�7�z�������^�� qt����%%�{)�U%m��g�箇
�{
�{
���M�A44��R�Q�פb):?�Ҏظ'��N8�) ���ŧ>�'2;3�9K�^�������dyi�W8%�%0���'���'�(+ 9{���@T@�t,�h��˺��c/��@��?g	��u��s
V�$k�|�zuy�:)���.�щ���C�N�������y`H_��&��Ø�Qz}��l!��._�2�	}��0؉&��Y�G�z(��{"���f*����1���#��Pk�n�
��x����Jw Q��4:��Ȇ!s֟���>fY�y��D�������FH�F��g���mv~x��ݸ�/J��g�R-�]����!d^ z����Ix���J�MA\'��:u�Ĳ�83!�o�R}�2��Z��Xb@� ,�� �s�)��3r��TG�E�Y�9A����1��0��Gd�!#`���L͜����d��MA拝�e�5�+<_�����g�]�Ku��٣Ͽ2%���ÿ.�,�����z��`�L3��T���VZ�c��^W���'����Z1�(�J�Aв��9:u:zkV�MN?t�HAFN�6��E�g9C=2��x�c`ȕ7�.�n k���g�t�&
�%�i�P���Q�X�e��r��i���ac�����I� ��pZu���E}�k�/�C>\��u���� ��֭���0� h�cf@�	Y#t\,\YRc��{��G�"�z��G�/j�p�z;w���q�[9�\î�)�}�:}��"ޫ9��tSĸ;V��
,LG�	�6��H@{ ,W� %9��ss��h�{U˭���/jlW��.��=z[���x�M�bw����^_�L�Q�	6~��8ݗ�b����W��#X���]�za�����S��e�l�rh�>�ez�1V�8�"GD�l?���Y#�oO�$���pU^Co�O�ݾ^��v�]Z�:n�Fp��D��<Ψ"�-�C�۶QV��g�Y��c
�Q�~���!���Ƙm���0�
{
2���1N�����RTE���?JA��@;3xB%u
�Ӂ����$WC@��#��=�|�u�����`��ٳgͩdR�T���1|��B�M2j�vT�iB�C�೾��jN��(����:�@�sp��d��>V��C� b&�e�r"�s:Md\���qF��c(ӡ,�GB�Y*%�e�]��3O��U�2���� ;����	��ܐ��F�d
���L�+�OJ�Rd��x�<�9��;|���N���Q�Y�5hC�^��E�b�G�)��@1r���x��g�ګr�-�ȑof@�u4�aS�!�I���	2lIo��.��	+j ���~����iN1����9Ƹt�a]���9����󣿡�A��e��|��������d��݃.6�(��a�1,�=�o}���'F�`H���ea�B駰%��Gd��<9'n������L2����Q|=�5Np�D��jY�>��|��'�?��{�u�ݩZ]�-��O��p���?��;����uvs3��ꛇ
���b���3�z͖��^{��STz~45j��UR��pX;2+�K>f'l��Yz8��Ӆs��� ���$�[ ��ɋ�L�qv��B��H�@�N�%�$��@�dW":	<l�V8��Mgݮ�B�i9p���=�������' �F� ���n,pD���PtǦj�3����ߨ���������w;�V4n��D<H��O�Y�f���o�0UD&��٘m��g�	�:�t��H١3��W��&�:�89F��H����&�#�5<5֘/D��.�37n�@���1'!eĿ���)�R��u���ef�b���}u��e�����_jFDY���h��N�؟��2���(֖�E_Ԩ�E���M��5�C�m2� ��juy�Q0�b�Z��3���Jf�~��I������r��8���o���W�w��c�&\��!��%p}Xs��Pg�urbTvՑ"���~σa�v����
��^�!�yq�s�a�Bv?�� ��M�[���j2?���%)� {���z�g�n���,�e�gQgrRj�������d��1𬖏��(�� Ɣ��5A��� 	�;�]/_f�����k�/O�O�rt��,��a��70YY	�H��H4�U^w�`��]�.<t�P�8N@����Y����0�ť+�i�L�b0�x���:��K�<���6&�>4Bu�z�${w�˻��^����vW���C���5_ *~f���y8T<(d�����ꗿ��[n��x�ìV��B �]�|�c�p�Y$  ���t���MGn�S
"�y�Vq�;���u$Ծ#�SQ'�LP6��Ϙ�3�g�r���x��7�7��yAʙsg	&��;�=Z�I����4��s�X��=935���6��J��~��;w��˅2AJ�0�=��R�HFW��h�p�o������z�m�;��5�Q�n���G�רG��ao�j�+!����ߵ�d�^9�lԀA!@vJ��03ZB�:�p��[N<�����P���gO�>ua�g7*�\C}M�������PQ��q���*����Æ�nĪ�mUd�=���R$���P<8� t�p@H�5݀2e�4V��*�@{*�����>�JD^ ��x�j��m��1��V�ſ��[�"ɭlm�*N)�klNj��؅�Cu�.#mO�v��a��S�Q��������v�K���q��(�u��NF:p��/��6�!��32��^f8F�_R�K��3�/�p�+��;̶�^��iK�V]�ۂ�u:ٺ�؞�Zva;��<u�Xm!y`62K#���ph�Z] Q#��b��I�2���߳�)ڏ$y]x�l��î���7$�Q��ѷ�vȋ���YX�pŀ���q&�%N��X�9.���ŠT�D��@+�
k����ll�r�#+(�b�ڈF��k}V�іN9��k%�WsLz!p�ȵ>��c����'���^�}>>�0�8�r�{z�h}��� �d�ڵ���<�kc�p�, M�7�O�5D��Yr�'-XP���+��q�AD��G|��b�� ӄ�wZ#{�g(z��&��t���_ަF�8h:�ۖ3R�3\���c� s�!��y��Q���Q�֣ߔ����ټQ~���25XP�A�s��c����B���VbΙs��O>���=��G?*��v��^M�-B]&t�����`{�ŀ�A�g��Φ����o����o�7��oʽ��O�T�6�ڃ�F�p�� �R�����+�?���8�J���%�O��}�eɏ������`pzjF�����z~��>+/.PW����n�$ՊQRe0�����=�R��$�K�G?�1�o~�w��_���'�b�|�f��l,@A�N���gv�Pc�jeh���r�=o�����3��+�?�<��lG`��5�z���c��?��������	��@~��������ɧ^��o�O�|�
�I�ܑ�vMC(ʈk����pN�w~$���.���[�x�A�Q[[.W]���sb�TLp�8qV��[o��.�د�
3u��Ϩ�~�(�f���d���|xJק��ΗC��sZ��G���>�!Y��G��^���*�2�=k^�D��v䖿���~鏿��}����?���G���돽�P���ICm۽.f(w%���D�S�����{A̋��]1�9>��Hr<0�66��[օv���imT��Q�y[5�4Je�az��h�HYF"ွ�YeH"#�Oƨ��zq?}�4;*��
b�'h+��j�J�i)aN�6&�@c!ѳ0�і����EW
�d$QAc�A�-ʨ�Ǧ_3D�!"
l`
a���ײ���`�'5��|y��=Fr�.��P��uQ@ɷ���Ҭ3�Bm�-���V�G�#TU���P0�{lRa4��(��3���!E��2l�O5:Z�A���'�ਲ��P�f��1�F�R95���Cn�$!�m�Ȝ��a�`�<1]��� p������G'aӷ{4�������5���r�ӟ��%�%�g����(���0�΁�� ��pYFbk4"8H���2��#��Q����a�}����95�u���4a�^:���];h4g�����<s�YA��r���^��QKNP`�UXkDK���EP�&]k����@�@w%3n8G�:�|>kk�7n2s�*���z�8�$^Z�G��C�K2���!;c(������r(VX��`���Fm��XnL�A ��5\�p.?��Uj()���g�)�'��K���=���k�`Vq3,�Dd�{MӜ�2)�;�����w���%�a����*�,�����K'x�Y<[[xdj9�]�+�g���? ����\��Z��O���<����!0��j��n*��������Buo}�rϛ�B0�>��zO%rc:z/1}�}�Ri%�x̜)�`� ��%�����<���~���O��'�H�Y�c�D������-�����Gy����ѷ.�u=);�g��뜔��b���M*nm�ʥ�|�#Gn��g�k_�[j8��]�k��-F��Y�q]�L ��:7�H�~m���}�/>�n�{��6���R./\�R�^s%�V#�YI�1��I��P*M����m��gN����/$��my����6
Q(��1��)
M�<�m=f5��-�,4h������G喛nd9�;�~���8=�̈qN�&�ȡ�/����#�{���o���r��	��W������[����%Q �{�;7�N)�����'Gx>K�ǠN�ֵ�6�ı�����6kh�  m�-�S�J���r�AF"�Nn�����Y������|����?��KO���+��׋,5c�j8^�^���窹�w����4�F<�Ol���wf�#�a�㺘�1����%q;Eu�5	�¬�VqE��$%Б>Em�ш�=��5b��9�~��@q��&�W�^�]��(�G����L�C|c����� v��8��u5f�ӍP��4�_���q=x����5jFt��U7�+q�����k��]� �����kpc�ۡ��f3��{x��"��!/ �0q)/f�-�6򛍴������Y����Pу1�����Ph[	'-3�����hP�ڔ]=_������^{]:n)�/�L�:7�S`F��!��5�����j􂰅�Ǩ�@��¹}�Z8>�*D�@.�s��/K*|ص���܈>c�lY��N!~�`����w��b@ �'���N����/�w����01�I���@a*�(Bh)��3��ci�*ObL�uLGY�	`�������${U�r`�@�]����`�G��k�y��>pL�f�h[���*-A�MC�9x�d�i\7�"P��>���\.� �>���ya)�?^}fY��H%`L����ۏ�{����׾,=��:P��:�NhWD���
@#������QS�DF�0�ʏ�A_�xQ����_���<��#�1 ����񡌠��߯�y��B�q�FY-��j�s^�����4hIʿ���9}�4�Xt�,�!`We��Fe�΍
��@>�E}���15:�N�c��Q������6ER�tw[$���2=�CJ�2��-dN��z͐�/j�e��i��/��ߕ��r\�����]��Gd]����̐��=��d��4ԡ�?�5r4�I�3j�g�2��啬[K�����:���Kt����]�ـ��1��曨�\����Aﰮl"��=)�]��G��#�~�N</���y�15)s�Sz�<q[j?��/�VE��1>�zkriiE����ʪ\^�̬ 4S j���edbd�ϻ�^�ځ={���C �Ҁz%��<����ƙH��(?�ޓ��0�KX�Ѽk�A7)���}&'S�㲰� �tϔ
��Ѐ<	_�ꎁ�|.��3c�rp�.m(!{����y��ɑ�����9�@=���Mt��E�7J�� J��G�D�ox��,,�O��Kο�ܷ���������f8�}��]��o����w"�C7�F�@Ə2q	vlM�~Q~�2*Nn��hp��.��3� ��Ed,7#�IE�ih�f� q��l�6�`��czXv��2�7�60�{�&C�:f� �62}hV�3�>�k&4�9��Tg;���~�X�6	S�Po�tL�@���nVdm����#r�*��Nz��n7lz.��5��������B��![�c�z@'�2�"��ԬH9:���@Dikmu��	�6�k��f�Jo��6B��ݮ��qvP�f� ;�i���������m�E yP��C K���MVy|+i�x���t!��R�6�:��S]QĴY�?���//�_�6�D-��@�����fBI�k!V�����q���(���G��esR�hU�ZO�%�U�� 9C��m�GY���0 �#&b33|��l>�t<���w�(;���R��>�+�t����ނ�����}N�����������+�:aV��\/�9pM�;���WLŶ���6�`Z������dl��c�ƙq���Φ[�-��ya&,l#gҪ_[�K��n!>�A�D)��)��:8T��,?��<�)}� ��[$�MO��Ը��p�JA&ED�Q	蜋C�\�y���Y8A6���B-���[[$��NOIF�%�ܸ�t��C�yp#
�E���.R�Y�|.C��9d���13�l�)wG��%��*������u�W.-��Һ�?s� �@��ׇ��o�A�������{�6#�$Wdl8��/�֥��6E�wx(�� X���8�{]�%�V�Q����r�)��t�kEfD ΉoK:��tZ���J-�(W��*"�R���M>��vbL��n}OV�W���&��i,6"S
�mZ1r�X���Z\����t�2/�z]c��R)lIF��QH�Q��&d��t����̴�޽�6��ag���.��L��H�F+7W�}N?FND�&�fdD���s���N�P"�)}�r�� Pf�'u�R
vJp�:�d5��6h��BY.qp?��F�B@�,Q�U#���@�xztHA[��V-q�5�t���wx$gc(��:���2~W`z_<u� #�d��	�t�V׷dbxh8?�<��Z��/�������������W�ݷm����A0����������闎����滻���z�Ou}3�!���[��������I���@�R�b���Ĉ����/����TNJ%�yKI&�(Y|uKn��y�[�&��t�>��,]�$/<�����NM�E�ɡ�5��.��F�Mm�l�$�Ȍ�s/0���e�`�|�@X�8��	F	-sH��� p�기(O=��FPg���
����!{�AD�Ͼ��Im����-�Ԣ<`����PF�9�
f�|?��(�/_e��e�H<�4]k�:Ia:��mH�A�d��U B�RW#^5�Vf�����78@���!�GJ �;�b��#ch������hJ��������Ĭ�vf!6�����"��C�Pc�	�~J�x:�>��~���0h+�T_�;�Iwl@!�̬F~҃�z@=�n���u=�$Uf��)d:9]�ֆ*(y [ ��S6��k�X+/,E�H{���P!���]�(�>H�C�����X��UL�Zm��ګ L����ۿ������ZK����1��w����gq-�e�p�-��� �m����Ix���$��!�u�� �#e���(2�P�T@��.�z*9�>�$�&d߮yٵsF��0���_�|���iu2Y � r-�O]#w�t!�A1tH�#H��^:� e����6��łM�N%Fd���sgYBy�7
��S�����g!:n(�A�]D-GmNG�y2��"�g�Mǁ�@y������q-`3=��r��������������r��vs�Ib&Z[w����ڦ��=�6F���m��� �y�!fo���l����&g����sӺNi遉�h���1��g�Q[�r�GB�����$��چ��q� ���p�Y�1���E���y�g�����*Z]Q�5>)7�'�~��;�#zM���0�������Vڒ͍�ɳ�A8ugt]n��v9�7�nK�h����ٿgN��f���t�\��Q�Y[�:�&��,�mw�M>T����om���-˫-ޥ�ob|�ϫ\ܐb�b�5�kP)��6�H�� ���-\�g#ؤb;f'�욛#zJ7����|�ۣ���}�|�6 ���	y˛���<�~���ɉ������7	X�����T2����k��{�O=�ұG�����3����?_=r��V{D���$�m�^�n�<{��̿�w���g޷��q����s�YO7g���Tmh��e�������v0��(��80	"��#�k�Mcܳu�`	uO��%?�2t��H�ԇ?�^ٯ�ԉ��/}E����H�Vu�@�������#7�D2�r4��O�]����@�q4���H_2���TF%�+�]�͚�rC;v\���SO=%�r˭��}��Qn<pH>���RE�S�c�)^�A���r�e��l6@��x�����8P�橠u��}F�� N����ö7�Z!���Z6�W@�
�C�w�lڠI�UE�'����#Ձ��S˔��P�I�"<�H� :�;I�,Mn?��&�
ѵ�pXծu[�؄(��� 2�^M��'1$6���1��S���bTH��%(�r}��:���1�<�����ćz�9඘�f����{1���a�F����I�`��8NKO�)?��n8)�׵4ȋ��+
`a��A��6j4Q��%�$l�c�7������mYǑ���*���ن���W����2+dU$�ڵ���\)�L�텝Y<$!���Vn�Z��J¡�1@s�����C�`����w��߀K�aa�$v���PH���
���jOi�c����}	o*ШZ�ڦF����2T��##���)ud�0׈�jNXCw%�`<�gn׎iS'��h$Xj���U
�5+[���v�5kE�M�(�ٞ9�@>�+��y���r���h@5�O��K�gp��"A.�P�Y��z��KsiE��A)�Q~N#S�<��7u_�RG�
���p?@-���e|d�\�V�Lǅr$�2D;$�w��I*�J��%�U����]
�Hy}Eױ"�jA�C?c��>�Z��I�$J� �vB��n�I)�͑\VA� [k����&����w�s-�QcN2J�bٽ�L���;o(��[n�AA�7V�(0����
��k��3 ��bA/��7�7'���&9�
�n�8�q�-�O����>�����`��28��1ϖ_ ՛o<"�J���1إV�������Y�&�aiМ����|F�p��П�����U��Gyj�NMC�4M^��̔>�"�
W�0d�Rqˌ#SۋY @�����8[�QR��Y���9�up�0���4�td*E�PQ�G�hng�Ә>w�p����z��W�g6�s����P5�HV�����^42�UkL�]�K�����ڨ��Pw��)Z�(H�q�a��S�Ϧ�8�OPQ�ģ	��h���@�Ь�(9g���#J�156*��$��ٹK.�[�?���-/��U1�r�W7�峟�3u�{�'''��Lp�z����#:�v	[HN.�1E&��R�owu�:z�}�G��1�g��3�կ~��.���'�ȓ?|B���E��/����7�EuRHC�L�AQDl��@EB}v)�\�1�~(�?W�6ȆG��$�����JPzB�~�]w����<��*�����6�I.,\$?��ɐ�a�:f�
��[�I�k=���;`�N��|�����8l��h�m�!	��6q52���3Yt���A��k:+��!�K͓�����a��A��E'�)�R'�����z:��=S��68dv�2�{��R���zp
�Zm\�7P<����>�]#�P	�]��OO� a� :JPF4
�R4��W�����U��W�����Q�~��u�u�jS��C��k�����Of8�J'�]���ֶ,���f��wJxO�,���}��d4({������Q��]���vE�x�"b�w�������r��mV֘M'�Z.hP�Ԡ!�r*�'.]^b sp�u�I��t�m�x�\{���j�&�YV�UW#^)H�^�F�@�|p�ny��eE�2�j ��5�U��v�dl8��&U����3ХDC[P�AT���#?%��|���\h�D��.NMA[yKZ�ѝ5n�0O�N��~��)"�r@��f���R#������d��G}][r�:hKƚ������h^֗.H�V"��B�%BQ�C
f굶�uj�@�ݒM�S8�b����];������v�����et#�e��h%~���xv��ô5u�pn�C��>}n��!�u�\]Q�PT���,!�Fv��)w�u�<����g�� f3������ ��q]+9�F��;���!X@�Ε$�ϭ
h����:.���`'Ρ�M�@��2��*01	du�j��obj�&���^g���� �r�|0�%Av �V�t���/����@�O���]�decCJ����
3{���h��X`n������P�`��{HfYփ�cwSDC��7�{�X=�ԶZ�͚�r�K=��k0K�ӑ^��4��s)?0I�fw�b�)�62΄S�tc�HC~���
T2j�[���j��R�n����P'$|A!��Fuȥ���)�����\.-\R#4DQ5t	A�gR7��g^�7����{����0��.�0.���	x�@�V���(~?5�Ac3~��_�o~��	�t��eu�4?���d���296���##���g�����l�9ƣ�3P�EFF���0�4���l3gC��3br�F,��� �3>>&�9|1Bn�:5�@�����I�\�6l, �(@�)8LL��HF�=k�l��O�FH�4�d~�:��]��9�ܳ�HhM&�%�g��p�wl���$���C�i�%�	3n��Yڼ��^B�������~)#R�)�����w(�a띵�ڄJ�Q8���1~/b�"�rK�Xp�Zi$B������<�])*�tT�����cт�L������ٽ�| �*�t/_��͂��9�
Ϥ�}�l�\GG�;`ŹF�5eY���/�����/�o1��"U� ���g'�x🥌���0��e����1a��b��:��w{�N2��S��硼�D���P~^+HȘ;G��6J�u)��r�F�9���%�{�Rh�c|��F����2���wݮ��)���t��,�m�a�SKoi��Y9��l�#��r��RޢS_8wZ���;$zǭ�>j�|�����?92-��t�:�Ei�3���ҏ��26���R�irZ^z�������i0�s��Y�-�~וM��)�������%��i�n8���def+o8���)dz6�V����*2:�P�>P�$����3�h�LdS��/�DXv��F��eҁ�m��lU��c�s"6�����T�sI�VMAA�%|D�F�&w�y��T��|~��Qt�plY���=�[�׮^���DiO[͆˲L�z���$g�Ϋ�ۅ��iWc�'t���#2�.�2� ���oH�+��ߧg����h��4S���A�n@�)��8m�7rU��F����zmйA����ͰF�5���Q`N��d(�uP�C��M��X[_���@p���>3�޶Lh���5��G�7�d�Q'�I���q��d*��4�>��=�S�H�2�GTr0����YO�CC	]imk��~N���̸���?���׽����E�$A�:�T;:�zc� �|��FŗՕMY�xE��;�Ag��#�KAJEZ�Qo�P�n�U�!x �R��̂��h$b�}Hԣ�h�4΄�ڙiP#�p��:�%�@�ub|���[�#y��?��}��TǤ8�k���� 0�l�*&z�( Рt�05�UD��G�Gp�M����f�i�˗��s/</ł���Q�P�%���� `�#�9�)���C9̳97hEFM��̲��!���D�I�Q���$tSjd�i�q�A^M�k��$�R�+����34�p3;� 3sԈ�e�ے��Y)�Qy#s{ef�~.^W�$�S�0�ϣ��p��=�G�M��	P���Ac��h�ߠֲyp��qMW%��}A)���=��a�Q�a:3�)�.�3AԊ�Y���������n�	s�Aȏ �ڷ^���,�\Wn	��*�23׃!�cI8U��W�h��R�c�!�9oɱ��dV	d��<���p� ����wm@�E|ײK��³�{S��s�d�=sND��:�Jѡy�^!�
������*��g)��c�5�̲g	�e�ע�4��;W.VdjrLΜ8f��D�%"p�@jt���[��O>.�xT��|p� �b�����\X�^3Bq:���166"��u��K2}��r����)��� YD�������Vg��+��9��F8��f �ww6�����癭]�z��$��"hU�j�p��� f�@�EK1� �ЍJ�5}�� �*� ��آ8فC7隖�%�%M�	���u�Wi����n*q9��E `p��p�]�PW�\��]`��I�}����d��qjq&~��)��f�f�����F'��2뤶*� �~��Zw�H���c��@�q��,>�+���k�������6>����F�g���1��m���&���C)��r] �����}�ry���h��{�T���^̄K�#`���C��9�~M}cIj�=�?��d@��±a� �ÖE��0Y�4`H�� ��x%����A��Ԗi����}��S�����#c��2w(/�����A�� #�R������~2� �m�D[冔թ��QAM����J2c��n��u��t��T��}H�x�A�xt(�x�������zv;(78�8��e����zV��b�Z�i` �dl@κ�EGg͎������ujDc)��p4<x+Bi$�Ψ�8�p87���r��(��4nE7E��<o5)�tuiEr�!�)A���ة׎�IF�d3���&�4�`AC7� �"�_(.0M��vr`� f��!2�s�Q��P�Y[���1������(/�Ǔ��EiT75j��H6/Y5�/����8qN�5*L����ufb��Ւ>�:ی1�iƜ֦�8�~�j@���z��6H�P��W��X���C��2	�z�.��,R�]Q�|}h� }��,�=:55�j蠥��)��D�)`2/��K�hr P��z=�K��o�1�5P�6,�jQ��DuN����N��>~��+�{2�k�����ɓg�4;��AlF��/�$�ÿ� �Z2�s���������\#��M�������/+]ו�߀	K=�r=�X��Bε�u�����b_c���P8�e
���3?�����֮�7�H����6$����8{ƥb��ڊ������%r�|�e���p-��Uu^)f�С��t&�gm8sh#!��y�C�n�<��Y�S���pA�z�����:�BV�H�֞���  @߿C���B���H���B�#3 _Bʾf�ãzv�N�TcܻX^�;��=������	������ @Pa5���֛tl�p ���h�e=���cW
�,ȵ�Zu	�P�9`�c)l���
��=g�l��Y@A4F���D����5�̐��FA�G�&j��� (S�*��\Z���9�1
�"eb�0F%�⾂62��� O?����UI5:|f l�wZ�:5]$��.���g�Ŗ�B�b3��lc�W*5�Kd��l��E�{@
�@�6��# ⇒�H��
&`_fg���yuyE��$���ɔ^��b��e���ڪ�왛�P٘�<�f'A�)��oD��W;���}���;�c<�#PN x�5`|H��&8�]U ���R2(H�c�\��d��[�Q7� �+J���l�	� �����D�v'	%����Zu%���H\�u*U���F��Vϻxe�L���i��ZЙ��O�:'
++���,fe�(D��]Qu>�z��lc��xvi@�P�tÊO�ݯ׻��#�M_Fݟ�����r��O;l,�� attt�?W�Չ����0��C�!T��065�H��0����H�|Vr�FE�=Y��rSA�xQߟ���"��¡As�^"slx�ۓr�p�Q-�!�s��7n�[�F��ѵ��n�NL�����*YK�-�D�7e��21�����g���3im��S��ճW��T�DV"����X�v씩�9qzAZ�d�4�D��U㉔-��h�tѹ���@�Y���Y	z#u�Ǡ~�5� ȡ�B�Q:�i�����4R��x��ؠkuW��LLR�.�Vwɹʯ6�L��u���r��N�mQ93b��:��%�EK7��Ih�^䡇��f�#t��I b��|�c�a#	�7�5�k��?�u�e�5��lCW��u�vî��;���觋^�}�SA���:��.�p�9�$�[:�lJ_���[C�p�Bx-���B*��>F�@!f.�Ib�j(�(�J��7����k��ƨQ�U�����V�HG �A�YF�؏q���κcf���EMkv���-S�=s�<�$�$�j������z��
���x�]i� ]��i
��{��}G>��A���^8��D�3��M<oHA�PnD�d��c4@hG`�Z'hH3�pm�
���:�=�HA�kekC^��2�l;6�
Yn��i����OMc,%Ae؍�����r�]r��I��8����0H�g ����f�)�����Q����*��M$�h :A͓:���a���Dc���4�#&A�5�h���U�ݻ�4�h����2Z��MZ�(�z:\,���M豃oXm{Q�KL��A�,�H@�
[�� ���i�uV��|��֤��C"5j%a�e@��(�ʒ���s'\V����e)C.7u�XuӚ0=�O�\տ{2:�Cr��x�<u�+�̾�5�Q喭��/ '��YA��Na&J��<@�9����Q&,�y̌Ǒ=i59�Y����Yy !0�絡���_Iř�gW�wјu�M8I`vZZ?�笯6�ݎ	#�C��Өn4X��"�tA��	^�+P��'�X��"�r��e���q����BQ�齵F�T�5��K��s�N��tA�׷��5ن�Cĭ��֨h��}r��C��z�20��	��rMΝ;'�/]��B��H$�x����w���s6($�m�/�|����ϚNK��$oC� ����~���fJ�u)JTn���mR7l� ӯ;��Z�����H�	#��MG����oݜ/�rl0�c<8�+Hۺ&���F������6�Y��Tu�P�������
R��VW)c])\�];F��{? o}�� �����{�hΓ���/�U���i=��%Y]:/�;����E�
�-�#;AU��R�� ��@��ߓmق;�0�)�$��}��I�=���Έ�Ԏ��|Bzj�2��-����em�
�c'������/s�����f����d�i.	F����];pZ��[�"J@	5�u5<pR0҈�@��O��b�޽4h�@d���D�Prã�6@�Q��8��W�o5pT�_�(�F�5��qJ��_nr��<&�˃N���6�p����CC�����j��K���	�ld��K�!���@U6?$ϯ�Ӊ�	aNN�X%��''gd߁C��3ϩ�-P�����1!���4�N���)F�p�W�\"�����"�@��|��7dmsK�Ø��"_��|��|V�LG�l���#>|u�
B�� ������e��s�Z2:>##c�l�G 25=kB�h�Ǽ�b�Lu�Y�G~2�#��S���tJjjW����}&�9�����='k�s�	�Ȁ�=Cl6 <�R����r�z��>����e~�^9w�4�u�xV���p�kE�vE9��9 tq�;yB
�C��Bj4��`!+n��N�Ò��ά�@��*IS��
�y�7��t���Y:���"�ūz�z>1X1���R?x�f�A�\VP����4(��^A�?���9#��㲴�I�q �R��)���ޓ��t����/�r8��lߗ\��$��]��a���+˜���)Pw�}�uxY�+k[�+r�=o&:��0�eK����/�-GJ*������FW��/u�,w���T������,U�����M��:VM �Ɉ�����@F���}�Q��Ĭ6���fٷ۝8�R��±S�x�DԦe2�>��M�̞��]s3��[����Trr�vf�|���Pm���%"I�럏���ޘ���������D#�P��e[��J]�¢,.[�ّf���n���#݌%�皁���o�`CR�bg(&���1���˃>�^�nMA�+��Ϝ9#O>��\Ѝ��<�f��}��(�Z�AZ��s����P1E=�0�x߾=��C����afU�&�ޟ}�<��w��ZgLQ����8tf�O��
�NKz�q���9�CU��s�w72�� � �ɵ�n�"o~Ӳ%؄�YD1���ݱC7��+E�&�'a;��k �	)St��NMuX*��lb4H�~C:���,�����
j�$!i��d4��TL1����7�ሜz吼r��o\�"j�{)�ե��r�H�Nf�̘l����3�Z���Νh`�"F�H*p˦�lQ�(�}�8׮V�褼!q)�=7�!w�|H�y<.�?�T52�Q����lU7)��Ό�{�غ(�����etb��/��ꃒ�"4t_�͡O��Z�6� m�2b��0TN#"*�C!�Dt�L�ݷo�'R�O(�C�e��z�Z�:�s�d��8+�~�Zk�����R0�m���m��;�Y�m�]���5�7��h�_������!X7@��:�Am��?!`	��U�+�w"��R�3 ���<��Kl���w|L1ֈ0RR�Q�>��nT��e�;.^Ҩ?���E�S�t��hv8���N�9E��ip�ёX���jx���;�geH�|�i$��B��=�3ej� J_:vL��F�U��j��� p|H]�͎3�Fx���.��,���� l��X�תrqqQ:ScT��b����Vז������*+�c�������aY��WV��¢��yeXC���	f�p
�H��37�A@�S�A���ɐ�AvYWM��r�����ά��]��M�/�ݩ��yv 5t
R+���Fi�6�5�Ѕm* �B�Jq=�	�1�^�`�$�� �jJ�Q`�v��#k���ŵ�e9������!��C�PLs�gYr�Qvh�����b�c/�w� '���b!MD�"�ݿ��q�I����
���w�-p5��Rc�c`˖՟-������A9`끯����9��F���ԙp����Y��\U{Z��_���"�{���Т�����
���9y��w�/|�m��R.^�%gO0��d�r�ݷ�{�����9Ƴ�cz�M`h�����z�� x(��9�@��-w)8�TDAj`|D�Ǐ'�M�Cg�QA�o-�NI���7���������Ǟ����Q����[8�J��R�r�/����D\���@4�2��H#�9:�9E�9��f��(tr|JfƧ���,S���DW�:��I�j
Z��&������)^K�P���ԉ���c�ɇ?�a�Q?m� �}��N�g&�������w�[(Fw��wɸF&��A�I����%!�]��=&j���`�e��=�(�N/�	�"Fġ���u�dkcK��y��A�����m{䝸,Cl}�;ߒ��י���T���%�;��9��A�?����C	G��/]xY֯ju�����Үd�y)�.KyuS��(����@FrI��az^���A[�ݮ�ų�8���y@�޺tp��0C���I�J��	}"G�I"j�fuU
K9��ZX���w�|�ޥ�"&��|�s�<(�|׃����sG��'4��A\�TT��y^|}�!���Rl���z�lGĹB۔c]��y�d�ú�=,8<<�S�M� d�n�_^�Lx3�!���&$o��I	��\s�}%���\_����=��۠[c@�ۓ���L���J����v	8o~���|]j(�KS!�	�6>!�'�8*�vf�ߵҗ	���J�k���ّ�Fzؕ�ç��@���9#���k˪cMX�DԜ��ZIj�9=��a'0�0��"�	]f(}�S�V,YW��Ȱ�Wd���#eu�$�_]ٔ�S�sM�gV��,F٣�{ �9��:��kˤ�4��Q;d(?%�QW*���Iu�%v�ml��Q�eZ?�����A7���K
4��w��{%�JI�]c :ddW���Ie�Rk�+�O�cy�\o��s����)~2mS���ؠt	�#��c�$,�^��W�~�da__Z���ّ�k����,��B��o9T�^\]�u��ܛ.����0��!�cck�QVA�$a��MT�D�j%S�{���Eٳs�0��Ξ=�fç���#�muuK�7�D��3��k�P���@�VW�sZ�!�����ԾP�L���UI�}����4Ot�ԁ�!��6�&���P�{~�
m88x�qɡ��F�X´T/)�)(�(jP<A�Q���h�D2��r傂?�< �!��-p7{5�ԠAmN�-ʯ�:��#&�#�䨽��D�gtAu����C�dq�G���/�p>#�)��;?�f�>���x��r˭��#���a<Wd���G���-N�V�xzM.]��Aت,\Y��/m����R�񛵠�<�V����v�#��/>X�I���
Tn]�,tj���"�����L�FS�uSқ�s,T�SĆz�nʢFũlZ�����ΚMd�c��Y/H_#R}����D�HWJU�ȩ��d,֢�g�SHPcp��ea.^\����&o|��2�)�����{����j�;�w)��MPְu��"V���%m)@�1��u�_01!	kS�S�b�"j��<�Xx����b� ���	D�4��6:�,-6�!$A���2�|���>CT�_:���:�d��ii/K"���K~[�&'��Q���ˢhL���C��cǖI�{|��ہ�8}NV�����4;2)[նlV6�ı�242'�l�ک���Y�3� ��L�N���Ƶ޵ɪ�t�bxkW.��s�uUd(�;n؏!N�������r�|�k_��G~�^������}O^x�\YZWÔ���z�\Y+�їO���"S�C�;��ZV����ߴ\L�����l|���UmȊ���Y����#��f�\��`@�*���\�h2#۵R�������+�gQ~����^X���)�~����n{��E}���}_����fi3S1Ȥ2B�5��g��������Dp�ګ��� �ܽ������s
�k�>��,�����2�q	8_ė���b�� ^nW��K��4K6H�c "������1yÝ�K*7Lm�Z�C���P�g	AS$��/ME(ͮi	�5�AɧK1G�і�x�8���ȨT5���6�8��RiL�3�8������T1��}�� "��3hq<|`/b�Mɞ�l'�C]+TX�(�Y��ڷ$�tE��@�s�����f��� J�鬍D	\d5G�i���C�#��Yz?�b��1T�H�M]� ��)	���s+�k1H1���g�pN� �P��A�AM�v�P��È�$���9D{��3g95���p%�$Z7;�x����q�O�5�:�Z�R�^��fd3�`����c]O�#��:�],������Į�Z�����tF�z?��:�Y?h@wI�_���/�v�X%Y?h\a���u�9,W��^]��S�J�3[
(3z���ע�AU}":i��G���]��YEha߷wUz��,�
2:7&�>(/?��٣�`l���9�쓒W�u�e�쌌��k 0;9�@�٩�ڗ�!D~LATb�N�=?/S��� y��t|����;~��n���/���?��i���
T�H9����;�꜈^��]L�k��U�T�$�SQА��.<"sԋ{P#ȤF0@��3��K#���"A�#�<"��Gy�Q 2:2i��PЬ�q�8�y#b!�P��Hd��\+����_~��M~�We0�mzz�L��ȱ@_gA1tG ��9I}��<�2�RS���4^	��lJp�� vw�O��ᘒ�cڹ �R# l�V����Z1^������2'(}am�9��E��vr�i�$�P�$G3�+�����*˗�P<KZ%�c���!Á*oV��~RV6����9SK[M8����O�;J� oNܑ7�p��YX�珝�7d4B���a�$�@�꾠=__��""#����14�'umj_y�|���ŋW���g䕗^��G��\Z�o�^9u�l./�}�dH#;(���x�/Xf��y��OJA#űٝ259,�՞��m�(V��8�d�k����8fCչ�H:�U]��BbE ����MuZ ��ڿw�:ɚ:�֫�r�n�}��3�N���&o��@ �2��a�M�+���u��(�l'T�h�-b-C}���.��
�s,�4�YVŀ	J�83���u�� ��>���xK�3�
f(��V�~s�$��8K���II�3��C�=_���F����@�� ��
�N��ϋ�Y&y�$ �G'eM��u���$�4�Z��*�v��+���QCA  "��?$_̈q�{Ү����`��es)�����\2H��qQN�@���@�B�_lP�~b|X槦��P���153�R�E���,�����v�r�P��� �fՉ������DF;�� l�ZYF�p&К��L��M�p}ã㲲�ίO��Sp�0�T�Z�Q�-��K�������]E�\af�@�в�r���I�㣺�)�_���<��ū��m�6a
P��:a�w�;�t\�$2Г�;�uAv+C��0��P^DkuW#�Q�*� ��H��n��f��u���g#�M�ª�!�n�Kh��dc����-��g߱������a$�3gϳ�SZ�k�P+J�ڋua]����ݦ���P��g�v���
~ ��C
4��V���ڊ,j`9��I��#���Q%(l�K^����V��BE�^j+������-w�䬕�@B��w�)�O��g/P ٭7��N6t`0e��(���}��7�q�����?�u�l��:*����dD�5=��᠞�ҍ����ظD;�@ێ�5jNx&�e������tI����6[#4��N�k_�:�OiԀ1R���]vi�N"�P\uUQ�9��A�ZE�4�廒&0�S��<��ìپ�}塞��6��vL�<��6������ ��@EX7e���[�cN�cz&��H��e۱E�@�F��x ��x�n�'0��XOF��l�����qo%�y\��{�WfU־W������ @$� ��(J"i�i�gf����eϜ����-ͱ%kD��`��A��HlM��}��ڷ���}y�qo|�����!��L�b���^����E܈�qIc�c��Uďt�Ѷ|8%�[TA�IU._9#�ν'R��4�� !�6F�!��[��ĖQ��x�z����g���j�"s��u)(8������f�i�4}N����n)B�S��c� p<OL=1B���=�8K�ͬ�^���i��5�����c�������*��6�mPo~����ɳg� ��y���(�L��L��3��������w���S��������tw��:������R0���e�����K�L�0�)�1�~��>�c�ހq�|6t�Xq\�`��e7:ٔ�w�P��iוi���`�6!�����b3zܕB}k�)G�Ծ�v&$ .��M��;:����v�7�Yd�ojL��=��27L�K�$%Np1� 4�	�L(޴�.��5C
jX��"���K�.�ޢϥB�+8`�$vK���d�5��ǞR��)�MH�����` �r�Mԝav<8���Yӛ����@��.]t�id�6�;y����ڮ�g�qV�}}����{,���"��@p��:a���!�3�������+�I����F�`���&;KP���-�XC؃�=�w�;.�����>�viL[�M��b�/@��ؔܿWΞ>%�L�,/�� ��k���� eJ>�����)I��D��g?;��z?GK�((�R��@
J��u%�����h�p�c������[nfk����o�׾�5�vU��q��.s
��|`�����G۷�g��ܳ_��h��رw�.R�m�+���{ŜąpZF�!�"l����<����'ԝ����?�����%g��Ѕl
�TW��s���q�C�����s�u�����﫽z��}c��$٭P�*�u�����O���]�7d�:ry���5���$X���l�[o9��G������e�/�ῠ
 ;h�xns��,���I/~J��]�jۊ
�q���or��]w�%���ٛ�['��y�s]^��>p��'��?y�<����Ψ�=8�D<*�;�R*)~��
aW�Kl����_�!�&[I����N��8[�ә����䕠���n�Y��e_�5y8,�sq������%���D?3e������w�Ò�G?��X��q��IN�R�3s�`��j D�� ҍ'�(p-JӷL8PV��XD����L<�݆�K'2,��KS��*��W]RT��vL���2>%�<W�o�]��P�,m4u-q?G�-�HUr�32w����u]��$#	���O����G����^i�3�"��{�u5V�u�C7G��"�6�j��ކ:��-2ړ��WʺFIC�V���ځ*����f@�)�fE��r���s�)@���#�t�C��{Q�P�	ֳY(�Usa�c��1ٴ_�{{d�$j����k����}GnU��*��{Q�[�ʰ�R�#؅�㬤F���
�Z��@7��"F{fhB�Q�&�F]��{�5 ��b#���e!�Ө��,�8�G,�}kZ+�/�X�k��\=�8�%�Tf��91AN�F6�em� 05�ƒ�,;"������Z'���?�o�"��5.O��x �י��:������d6�����{���ŏ0#�?=}���e��=w�+���f�X�|Q��B�C�(���ݧ6�8�stԁk ~�͇����=��+�ȕ+W�~�V��Ո~M�Q�����c���N�g�ق�AƝw�%{����=w���.F�t�O$�D�b5O��_���nm�� (p��"�jx�On��6y��wdQ�XC�� �� ��ү~. )�o;�G308*=�Q���%� �0���5*���_����ߕ�o�G�p�����B��L]���`�0��>�{8o�u�&�(#�g�����o�/~���O�v�"�k[� 7�����M�$Z�UD�Ȁ����r��e���?/����O����rdg��z:ũ��K4	PĮ0�!���,?~�9��G?,��_��������t�z|뜳�S�bY��#�� ���B9�����A������_�?��{�l4�\ZC
�q����A��� ���c++
�>�˿"����Ap{�:�i�yt1C��Rp��xt�3z�
��\����R�W�%	É�1 ߲A�xL�r����K���P�;#�.\fFnlr�Ā�n+���袜�|U^;qN}�exl����|����Ю)w
�&%�ϣ�[��ܱ�H뉏�C���_~d�K�X���.�|��1u��"�q2pPCH��ͦ�Hڗ
y �l���;�q�ѐ}�!���qT
����:5p�h5�b�'�+�Wk�� �A�4<�>�s���o�}��MYe�Z�F#uӈ�Q����F�2I��*����<`����:nB��)1O��tRP�T�;n�C� 't�dՉ �B���Gn�+�h�)B¹R�OPwE��>vL�=��ɢ���9��+�nU�)��6� <� �_�z��r��2=?'+j8���<����2���d�$�V�_[���/J�ZDfo��U��r��^y�����ʡ�a�@b�)��gD�-���٪��
%\�ܒ�.\�d�h��M=
Z*o�e?#+���(U�݁��j_���P/�����S <>1,o���;t�L�I��5�t�l�s��J-N�� Cγa'd�b�,�Y��RC��~�Y#(d�E�/��,c`�;I�P��<���aG���i�{����>��\�N��&Y��ee�N���E�g؝&V�2Yu+s�\
M�T��B]��V�OL��>�LH�-v�2�v}�0訑�9F��c���-���'g�2�e��� ���&N�dϝ9+��{�}\���:q����A5O��,?�x8�vC�;��F�C8�}�n��}FvF��W�X.\��R��8k>˦��t@�yk�D������T8�_��g������v��-Tg�T�ׁ���4���� 2�_����[n�����)�sE�&'$���9!Ȇ{P��#K0���@����s�H�EI:t���q9s����"b�� ,,��4��]���ÍF���ba��>͜3��ŋ���ޔ��zC�y�-v��)�#����Wi�HAM�~�=q��+)��A'��܌�@����m۶��E�8�	e��6 �bm���|+�8t�}���ӧ`������y8�w 8��! �5����L�^V�#�5�{�T������������]�����a��~�A4�@�"]P{;����?�}���Ik�����B@���r�`@�S����֩#������{��z���7��ڿ�|F��v��\\��e��c�C����$�^[\��}S�6��@�}-����}�VT�M_���/��'Ѷ��?%y饟��[���>�����|dV�	^7����s�B��Hn��`D ����a���D���a�cX�\����/��BUG������ޗ߬ۛ����s�y���� [�ah�����h��=�Z/-�b�.�z@q�v�0�7l�������#3:~���C�R�~ؖC7Ǆ{��"���� c=�7������{�|��3�e`�#���ʃ����A�ȋY�д)<�� �����)+D�#����?x@�TCv��iYY�����MnzL�Nl�&�#$�":���
�>��sb�1u*�d�F_�r�A� Z k��Q8�&��\j�qc���s�[]=��e�	��H����gN��o۾�zq-�5��I�FЁ��k��V6�8+3�eYW��Ո")�L\�jE5�y��A٨n��n� >M!F
�W��Aг(){֎��<�6�3��v��[��}�1���x}{p{�`�\�7t䴻y��yټF�?
�d�\��� >�ϻ����eAVC���2��:BwN�u�
6/�yD4��uL���&�G��}½�-'Rc�(FPD}�4�k����̃�����o��������ףN?��� �#�Xsf���������>%�_��oP823�Qt�C����R/f吤�� -��T�>��7����O}�Q����L@.������`���%%7���{��:~������|�����O~�%|�Zzݙ�me��v��sD��p��;C�煗^�W_�{��4��j��3�����S�IP�,D���^E� �+Ȭ���,�2A~{Q<� F��,���W^3{��j�z���J'���!y=,a���c_�L���P�e�:JY�<�<C��A�� �� Y'����_���W���,��y������|�A�pQ�c�h�M��`����;y�LOO�8?-m�%�1�|��I}�i�7<�M� , ��e6!��Ac	�G�,p��<|��>o�U�]���@�����o�j�A4l,�ÿ��Q�^���Y��9}��.�O�P��q�ª��-['i��i�23#o�s\m�}��C�����$w��|��Ɏ�a�))o��/�=v�PX}������ eZ��^7�L��դ�d^��}a�b�,1�9�m�hQ��|ڤ��i ��7�h�1 �6��w�A
�#c�M����h[��6ZFj�r��W�lN�v.��ӧ��>u�L��F��.J�zk����u#իMւ#Ea�/$�[6��m�QE|G(t$['Yn���y�s���5E�D�^��4�Ҍ��1"���a7�H`����ᰶ�1�M��P��%�T�h�G�	N�=�_������G�����?�+w�s�?��ɨ�ʀ�[�����19q�tm�bD��e�Z�{��(s��)��,�s��,���KlaN$<�� �aHR��&��H�7uM���\�֡5����gnuA>��G�CZ�A0�5�k
`�����G�v�(#@C�%1ކ�2��
%Vf�6��]�iC�c��� �L63h��i;7|P�h�\����M*n{F��j�?�^˿!�%�E�-�1㮔�9��W��	֘L�:�8/n��&�w�)�v�|�^r��o�0�.��"�
����XC��CN��,���n���fҼ7D�O=��<�쳒U�[e��N0;99I���jD�<�h���`�s�,ݾ��;4�8���G���p����e6�$}�]j�<����]p�o�����?�!#�=�E���3�{��2���u \�z�]��"������k�,��=E�B|^b4����!���K��*`�X?����tO�4��u�eq�>��6px�f���d��N>���8}7Z!�JX�Xm2:.�p��Y�Ϯ�6��)�yQ���
�,���%zqm��&�kf(�V�؆���R'�u�Tf+5:��>(�l :Q����0x, KX+��	l�@�Q(���I�{u�6�;�=	X�Af�=�*��R�v�?��N�;Y6��Q������p��,�@S8�a�#_�c �+9W�%������z��� h,�g�[�����D)��ߒ�����<m�ﲴ ז��B	�(s�A��Ĺ��y1鈈\�����g�X6�粙o�7���ڏ������_��+�O���@��X��E�Y�(�3�D��D��h;R�E��!h���Ø��@��"k�8D�B�$,�ŋ�뿈O�����T��A�F�x4���*`x r�����-����r���g��Zi����L��6E�e�[��*#PF�׊��2ѷv��Qr��t��PQ� �f-�>���ihA�C��x��s�p
s�YΪ�+�#O7$�����7��$��WY�G�?X�0��b����'����a�`A�^��U^FO�)����U�,��0/�� ��Q�: c��0uL�W*���,������X��L0 7Ƃ�����`����՜�vS����	�����g����9�!r�^���1EeK˻A{V�K��x��oapa"J��ÌN-p���Z1����!��r��=�EҞ�,�6!�w��v9��,_�m��͒��kw ��;7&�o���y��M�Z<�(�5���5/"�}��gC��D��u+�5*�>�	��#���M�E�y��1�g+��	�mr�:G��.J��4E�I#�A*��'��&uL	֨凂�F2I0�N:�[3˘F��N:��c��6��78!q#/P����҆�@�e��C+,�t�7�6!��y�Ta�6�Cp����y|��^�IвQ /� ���6W����y:��m@�ɱ!�=t��g1.oq�;;A��+�7y+p^�*�,p8k�s�Q�7���2�}�M+̀{G����L:�{�pn()c,A��d��L���H�f�6 ��
�gCq��������� ��������L�	�<�fwDB7�/J�3B]A�k� l�o���)���i�>�d��0�(j�YQJFI%bb�`+�G *�F����W�� *����a�X_9��y0f�I��zòK /������?e������؄���þ�8A��Yl���ɇ�L�V�#�"��ӧ���K�eb�e�~��� X�+ϟ�z �GL�qlx��v�
���۫Kk���@��ҽ���pQ������t���s�r�z7�,8G�K�� ��j%�^ʝ�����G���׿���t�����~��5�S���;��r�7��M����H!ҋx�fF�����ÈTҤ���Y>l96Cb�ލ�w�קέA:���&]����h-���g�q8������x_�T"�F)D�|�5��u��7q%dIh�]G^4�m��1򺔾[/�#3�M�v��9y��O#������ٽ��(G��ګ2;?g�n���{���ȹ>ӏML��m^�Z�絜{�С�t������N0B�#}��������F�x&{o��ai��2�Q3�������Z�e���}�4�7(_�x���u-N��[6��t���&�d���|�u9s�>�і���P���(��\X[f�_����}{��	��"3��ك���b�Mq�-�����a�F-B!?*�03�<ߨ[��3e�m7��=��dS���{�e]�d:fUP6hm���A�)d< :7={#�:�ο��qz  y�IDAT- �C���,Y�!vh�ޫ��w��Ϡ�J(Ї ��r�jtr ��e٠���l�����ѣG9���$X�P7��V8��U�0�/�{��z��qp����<��s2?;'����q�\���u���7������Ʃ@��j�ď���<��d��}��#��`����D�\�v����z�j�g�cC�(�|���裏���Y��!p �.� �BZpx���q8��쭷ޒ;�S>���L�f��KPi�3b	�d�p�m)@XZ626(���|E�~�y�[Zf��j�7�$���4~����r�*-��*���Z(J�s�vۭ�?!{v���g�
�g����2q���g늵�e�'~�$��?���r��w��9�Zf9	�8����� ǆ��
[��rۖa�:=���l~��'?m�\w֊?�D)%M;e��%���D�K�8Hw�q��acq]\��$��Gm���B����U�ro���˖!�wߑ���q��w������M�6m�M́�z=�m��>=�(�����TS�ŕe�R�h��L�	L��*mT)n�MT����x��[�{CSk��O�.�꺷sE���Y���b:2��q4�4-+�7�}�V��OON�?��O<����O`Nn����f~�k��3 Fҵ� �
!1��8���I̙G"~硵S�m��qE,�
:)S�~۵|+����¼��"h�{����Ⱥ��)c6���Ƶs�N��ny�� ��{��:���i@� ,,����s��}@ŗNf�z!D�7����0n��{D��!���n�ݐ����g��|qÈ�������!#d���J,�@@�<���*6i�1�>��e'�KE�H&�֨v͡��G���Fq9ɭ-�D���p~o;��o�TB���#֡ͨmƘ�I��,KĞ)D=l2j�R���ڂ9_�|Q�]��Ӄ+聄Bh¥�gթa� @�4|'Z9{R1����u��0�9F�v\dyaU�F��n�&V5b�'��D���
��}��Y	++Ra�INǨ��F�Ɩ��� 6]km,a��/O_SP�<,�eN�R��$��4bG~�l�6g�)�z�r}����$��;��;�L�#VV����j�ۦ��G��lߺ��*<�޾Q˒�@,��C#e tBg&0v�;�GG��O����h9�3A7]̏�{ *̘0�)nBh�5(gvg�!%�÷0"��9r/�����ueE�r
M���ŷ��G�����#Rvn�F���	���A �8PX��
'��d�`�x}�� E����[o��m��ܺ�ڳ��Ź�E�)8fi5�)�6�	�=��YPG#.X�R�|�m���>��rם���L
�x΋iXG2�fM�2{��0�
{ѲI�P�ݺm���n����c��g�`��b/�% #E���{���2�BeWL���ɗ��%���[ߔ��%�>E�T�Y9�� @���\'�88\r�k�o�>���>���3��~�[/����p�4�7�WԦIZv���2u��vS�-�_��8|����T���
�1������v��T u ���`�@k�.�G}������'����7l^�glYI��t�&)�ke�r<=�L��}�����/����ɟ��s��/��/��w�qP*���y/�E��e!���x7f|�ٟ��|���)'N�����{YY[U[���<8]
X�u�~9l�=�9#��,ʽzH��~�G�G���<h�)`��Y��t9��n%HJ��Z��w�p���� 忺����������3�hJ���p�7-���1��5i�V��ű��+{�3�Ġ���m��3��]���i?����ݠ4ڙv�m5���=�|���H@����*�yjv�:qN_�3 Yf���l�NjQ�l3*�6Ӗ4.��i,��j����W^�����ks���?�2��R�/_�g_|�yVw�$I�ac��c����w3�p	rW�F�w�u��޾M�]�fgȌ9ã��9�4b{wo�͋��dRQYW04?wMV���!�V�*�Y�q�� �;R�脂�cH�Ώd�R���y=\��QX����Z61��� '�*~&�[�g�p*�5e3)%�|��W�t�0��]I�_��Qm�ϡ��(c��)5,qΡ���Ȑ�v�f��95D�0te/��_��0�0|��J~^g�z(���\ܔ����`o1�Bg[[+���63sn>�uw@%�Qk	��
�i���,�j�>� e׎��F��o0����0�
�MQ�n��J�LJH�ozM8��>�!v���G?�׏�4�@蛠=��$�k�m���bt�n�E����������[tF�>��<��'d%��y&!20g��c��`��Z'8�Z��t�'���'��'�
ľ��o0��h�N�	dML~�3&�JL���a�XA�]w����ߗ�-"_�뿖��~G#ЈTu��@>&|U�t`(��\�h������^z�%������Vy�������>;�HȆ�c��~ۻ���iviE9�&$X�����?�)������~���D1Cdt]9]&��umq����XB�iD�����=ǔ�C����U8Ȫ�/���m�q���Y�[][�Y��DZ�=���/��/�@��9@�愈�vq-�Mt�@�B"&� �1?�������K]����|�p�x�h@ ��Q�8KMޏ�Ԣ�@��{���788l�!�V�&�s6J��G�N�M	�C�%���o<&_��o����Ф��0[������NP:Cr-@����D0j����/����������ō����(�" �c.�>�Uu�RA�D�.������o۪v|D"����yjŐ�N�e\�x#n��G�ҺtQ]rqi��϶����۞�ʯ=�,7�uc����h��
N<�0�=Q%N�u2�`�D�\��osT�C��H>�F�Bd�M'^�̞x��?���di��n!�J���n� �m�P���]l�h�D%�~��͔�{LCUd��	Qb$�Tg�8�Ydpϊ��|��Mh�a�*�� &?MNNh\dn�]�A��`B��5MS$#��XtBVC�&��.�]*��R���Jӫ��O���4�㐾Ŕ��j�&�A�D��D
�g�F�j$��l�{�
�%ٷ{g���)]�S�%��D�۲&Q�D���`~Q\����趁�e� u]J�:�K|����(Nۤ�7������e{�U%asj|��=9}f?~�G
�9}v�z����tF �!RD���v��^+�:J��ge�b�m����Ǟev/s�4K
Ug�}�-7�uʑ�h�����b ����&q��:F���#�E6�I��pÕ�����7�(`,��ӑ���[o=,��=.o���7�X"7H�p�k@u3b��^�0Z�c�50dԓ'����ޱ�]f���2���WS�0��d����С��-�l�U�n8�l���ӟȕ�3Lۣ���1��Q� ���b+,a!�����6Ν�g��������{r��	N��6F(�E�������	��bt ?o�����%�ڲU~���0�8�!�^�z��	�\jrx�!0�E����1�H���O򺯾z�AJ.�r �6ԡ �Pg�=s��"x�&	(	A���~����v���E"�밤�f[z�2F��l��9[\�k�<��ӗ9��@�,>l0�>�yB('�3��F���[�����U�(���}]�(1�9��9�����z��z�E���nYhd��P� ����_gy@eY"p^�5���g��#���/�4�&ˇ,�+B&jyq��]��Yt����
62,��w	��)r��Z1��d(��`�q��7�e#�	�L��!�Y��s�<�Q-h�H���<�� f�K  ��ȸ8� p��+4H`��X=�� �b�$4upsȑ[�L����~PX#}�g���u2؛�M`�Zȝ�<����y����������n0���.��{�R1B$� 4BV�G��.0�	�����ĥ���a������uh��\��Mv2G�;��7)�Sa:����זh�ڡ��Y{j�x�6��ҫ0���`Ssܸ�Gs]P&�ږ޷9p����@�׻i�u�H������#�*�Ю��B*��:�#ɐ<�ȃߴo��p�/5ڤۥ38�v�c�q���l*�Q��ؤ��������� 21���F�ӏ>"����^T�s��I:����t��޵]�����yy��dz~U.O�a�x.}}i��	�� ��;�(=�1�>�l�F�}ѯq�x��| ;w�!x����BwWZ\�#-�����T����K
��eb�V�z��8w���������i�d|l���Bn�� k�{���K]�]��2f�� �ܹ��ݕ�f��Y'��`�aL"䞯��iw鸬�f+��dY6u��ōj��%�\B���}���s�D��>���,�R��N-8�r�h%-��8OU�4�:-�i �`F�ّ�����О���v6��н64(K��
�W�ܝβ,ؓ�eYomi�ep# x��C�N�S��1���'Ml��9�����7��c���|���x%x1ӡkΆkqo�l[��g[:��z���Ȩ,���=�}�5:>���0)�,��g�S�-d��t����Nah\k;mv���nX���!u.��$�y��c&�����ɤ(��-(���߁,����A=j��6"��w�f�'�I��i7])ɦ�uB��ݲ��qc�&��R6�� J�̏3���\ �T2���A�Y�x��� C���{�"wV �=�G+��ש�[���Ȁ�,�^�-�h�ǳ��6�V��6gK�\�2���.��'�6d��̠��mldȕ+�X��x�xDfl�gF��g������t�E���~�#POH��uj���%=#h5G0411�����w��*\�D�⢢��I��CɲK�ʛ�-���U�m����yн[Y�v���	� @�wH�����+���Ɖ][�~�ӏ|����C��p���&�&es&k�6w�4X��!�$nCcSvţ�2�1�ct�ͦ9m�m _vapN�����#�yd�o��f{��˃M.���6����.
�Q{���<���,�Ex�uD,cQK��4�He~~ϥ	�"N�4'E,��"ih6��|X���!���Iٵ{���/[k���d�:H�{q�0'��^0:C���D�v�jN���@3uP]]	����	Y���aKKR}q)��9{�����.�w��m����{������T�K�3<$w|�3rˡú&q�'�zVf�4b�8ν&	�ܺ����z��� bBIh�FD ��CZ������پa)/�H]#����K�3r�2���K���a����
oU�'J98̓ȯ|��r��w��ʚ������o����\�.arP#�n�b��`
�81�-/M��1s������^����F����E�??3}�ľ �:�\'�8�9��g�\�ڈv����	�L¤�J=�&�ӷ��|�]��n�<���"p�nFA�g����1�4�8��e	��6ޞn(v���l� +E��'n��̲��Eh��K�!Xب#H�ѹU㼛ެ�rB���,(|<���,�ŚwȷХ�s	fw*��"�)���	u��.U������t��Ԙ:��4fu%�Bi���\@�so�&ha�L�dOD��EG�4HP���l��
�2��1���%�R��kA��Q�+��F�;{�GO	R�z#�.:��x��|D�@#�T���B}~x�)��>;� (lH�v�Mm�	���vU��B���`D�����" ��f�ZM�D�=v~!U��h�� E�_�!����V��托���#�e�) �l����4��V3��$�!NCbϢ��S��\2 �ra�D�d҄:#z�U̵A��W0B���-��~(a�������3  .c��]�=/n��g�(iӲ�3Ğ!ȯV����P=YO:��m.י��ӣ�Jz|f���j�/S��0( `G��@�	Y��dԈ��yv��(8�yn���7�x�X�w�_b6.5I�R�B�Ha��^�o���9��/<��7����7��s���E�����N'3��f�LF����#���9Yn�4�u��Jt-�q	��뮰�������Kq���=�Q�0��_;m�$�5�B��G�0�ſ��/BMԃ��D*����L�Y_L�����t�P�@�g���"z��pm���o���l��<@��F���]�(��JN>��#r��}r���q�������^T��X���:i��ICL�g�Bl��Trz����U�Ԙ>������
�,�$��g������{�;�<l�����ru~Y��n=$U��"[w한�wU?GG�3=����Nn�!a���R�04�U�f�I+_���i��ko�%�s�#m�H�AI����R�"S�X�������ȑ;�H����/��}��~��W�9�ndr��X ���w�7�9����~��Ɯ2���m�"i!˕͖� �e�:*�R�,ںN��ѷ7������`h꥜!�EX�l�9ۼ'�v��s_�Ϫ�k�ޜ�,�ơ�0��>�gQgM�7&˦�	FYA�*A����A'�E��,��H�#�����hV�9 �׼8=M�vJ���&GP�g5>6� =A���rN�:\B�,i�T6�wWI�	�D��'F%�P�
0Xv���k�{����Rq�ae�ޣ�\�`���9ԓ��A�=I�ٹi�v'+�	\��L �����~�k��ד��
���ʒ���k4�У���� #�rMV45�F��f3q<����ccĄc>^�X��y�l�Ӏ��= (�e�aojm���۴g�?���݁��4;-����&���g�}�[/�WH�6��ϳ�'�����C�F5�r� ��	Y�3�&��ΤHRFkq�� ���"Q�6�(A000(}��,�}�J��
 	��?��1${���k��j����BV���u)a_��u@��7�ڌ�Y!8ͯ,�k�W��{��=-���4r,	к��9��C <؟�����2��XA��Uz��H����;b����p?S�S�9�׌?�!�qó�@0���c�`���^�"4\D:/5��Y�(�*�<��AШ�7�vM�����
R���1�
T��"�$޵iO�a�[�j��лFN�/^�`�G�bz���Pq,���ίh$�̀��R�U��m�h�1
��]N��xwW���m�f�����{���C��*BZ����Ro�7�V7�&E��bjH�b�*�KT����V����͎�%z�W���p��4��>�DԸ)O>���a���8����SD�S�4�=�F�ARaS�b�}� ���du��~��Aif@�pl��rN�z�ܼ�3��\�,�����LL�Q��ʕ9ٺu\b6:I��S��{Z�-J|d�l�uP�t6P��k1B��6h�Nx&�p���4B�����FA�_�z��-.��-�c�WA�����o�6hY���奂�>��l�/z��w�ĥ��z�2:�E#���������m�NT�R��걬OC�$��-:��\ӵ!�Ə� @9��9t��v6�:+B�@�Ϗ���W�	�Bk���(�{��'�o�t|<���)5[1��Tg���@#O�4Z� �PJ�j�j�ׯ��W{���LG6ۥ�4��+d����{�Є����շ�����7y�}��(�&�a�m �I��WV��Q�(������nuHٞ4���t?��V݋����Is
^�l��U�
� ����-��.��ꊡ�j�PÍE�QSP�tq݃a���B��>�\�����U:p2����z;��
�S�]�2�/rם�q,/�&��^��~��-��*�&t�c�2�}�8iݿ��h��Ή��&'��ɓ�u���V�\�sR�6X��׫;yw�T`R2�W��9�c$M�Ĉ��-�m��:�(��P?JwI%�4�Y��l�r��uI�=T�;� �Ae6�Uvɵ�>`+��{AR�0^�����aLwO�uP�H��S���A�}�������:
x5(��`�W�7(�����HJF�%��$8G�Ef��'�Ə�g_o�L���>I+CI��xVU�,�[��~�8S 0fkt;�� �B��dA��&V�-Ξ3�'<C�� @Q�W,��y�lup4X���U(z��'�©��[�)��t�d@�k�W��������}��u��ۢO�4C��Z�Ҡ,�B��l��b��G��s���nxF��w�$��9a[��2hw��(!LK�g�%����=�vx�>f3V�hdׁ�^ٻw#�re����s��M^J�,���˾�,����d�´�����w��O�9��0!���e�´\:/����.�	�8�l^`����uF�st����5"	LLj��1rzt#w;�B\�P6��O��$��jh��e�*I���wD	� �Tk�4���B�,�42*@[��ѮP���t&��)�	��OQ����o���U�������g$D���K��Yȕe�X�HZ��6��������!֥`jC�#"�m;��g�r�b�!��/�7���(Sc29>�.0}�>��`j^����W����="QY�	�� �>|Pư:h倫cf�c� 4`
wĳ�����:��27/kk9��m@U�[���.�� WRڻ�#l�.���߾k9����q����u ���ｿ���=-;^`t�uo ,p�2���j���!��>��&��G?(?x�兩��];������dM|QovU��-�fu�����'�c����Cfk~�WEANV�<��>��ٵ��S�����Y���0O�b���n�T�����rr�1���a����y��#�.�'�����6�G�+��Џ�	�2�!�/z�
D1,O#�ޞ���ܯAJV��s?~F��GX��reZ?k�l(@����f��m�K1�� H��*��n��?��ߑ|�q���A�t��I=G5<=�&�Ydi�~(k�4A9d@�R��G ��K~�������LA!�!?}��[���6��W+��̠�s�s Zע���Y�e�=�o�r�ckj��@G� �*��lX�Jk�,K1�2u�R�YU{Q.�dT�4r:���N�7S[�� ex k]Z%t�E$��!��H��)��SY7��L�h��?��B��M�:.�l9�|�G�/�R
!����g�`�� 8�H��J�NUX�Y�ƫ���e��]�b�>ˡq���qƔ�'�x�o`��^d�Qr�yB��������;���� u��ПEy)�j���jM�j$A�jbd�g@�\�@ϰI�ט�όrh,�M��yC
h���� XAW�L��X~
��'_��{a����=���*�B�_$�L�����f� M����5u�,'�Q����^�m���RtG7���N�q(d��� 2g�Ï�nI;��j���_��o`A:e)���8,`�C��e�b�G:)�9�����ڴ�u�S��$^(@�@�g�)�i1����+����BW���$E�(<�a�Q�&���~5j��ȡC7Sz{na��R�U��7��͈�n:*�"SA�G�)��hd:�c�~��Е��Y0�o��ʬ?��fݺ�:w���఼|�YR's��}������:x��MJC�
��q����-�l��1� ���i ֵBI��j��BnI��E�	Fo kp�(�\�t��L�
@�ۀ
�FN4�
j�\�"��,/��m9v�M��n��p���Z�\d��ď�G��*i�;�I����4eS����XOd�HbnwZ�m�a�8)��ˤ��c}�=���x�v��A>@��5�Z����M�nm60d�].�F�Ƅj��V�Y.p���  �k��h����&��YJs���p���ȡ�q��9j��P������Q���l��Jy��{e��q�t�Lm�/���̙S����q�=���FQ" \r	PT��~:�ː���{o��[{erlX�a\��>����3R<��{���M��%�ٰ6Xr������
��������^9�NЦ�3��A�+���k@�sin���~Pb�tb�{��7#7��*c�t�2@�]*�ШI��r��3��c��\�Vlў ��!m��-�5>2��&F�5����|���+������x cȂ�dItI%�v 虊/��xG�'�=C��̈�{%�ʳ�?X?D���T+��P�Z��~��{��J���r�9u�u���9�e4$���hk���S�������)���l�Ν���k���� `�Y!�V�mV��&\	�'/�N3�vpa T@~a�=�c�=<W˞{���~�)�zm��3�K�9 x�bG�- J?�,d.���5Df�+Ў��]R�N<�p�S�TMLTL3݅�(`&�j1�.��*u��앺���+W���|��� �����پ�|Q���W��#�^s�`t��Kt'"�̍Ԫ���������_;p�.��׍��1��{��nvf�X����	��-uuǘ=@�d�e��F��8j�uF�;wm���&��p3V��U�_x}F�	������T���̐��ǯ~�s265���91�6��$ps*ڳ&0�Q%>f�4c���&�6ڠ������Q�q�<''��>��E�]���y�$�>��	�A�A� ���#T�����2%���@@G"1"q�����B��sUM#kxܜ��HvP�aX�K���y�F�'z0+�Ja��zQ��JJ��dZAT�'G�o�������28�Sz�����}RlƤU��Du����#�เ������� `ܧ����ئot�Ll[�����s
fV��h�X�1�2 2=�x��Iԃa\s3
��y�[�o>)U}�޾	ٳ���"�+T�������&`^ƶ�+��Cv��"����DMy&U�����۩���2Z�[A[tͲ&^[ 0� ���=p)�vyѴ��m�1F��BH����󳃬�w�H���*�X�<l|v��Bm�{^���`�ܪ x�F�[�<�<1-k+�rmzZzR��}��0� X .�Q�c�g:�V�$�]�Ãr�m��_����m�RE{���+}_�Z(�����*��@�G"-:D��z�\����޴F�}r��Uv�����O_���Id�{ �����Oؾ�<�Og�b�Ȯ�{9廨{*���8ڗ!|��=�3�@��Lh��bľ��&8=s�kAw\��ʲ�=�g�N}���S��:���]����}~��u�
,_D8"�۽
��Қ��r������;o�+��_c{)�A��+ \��W����m+,���]�7�5'�������p�*�������h�l���0�j��wKF����7Z]Zd�L�Z'p�j��!nhP1�m�]bO��w5�<���P�5�Jw�*�Zg$pl���VeW�܅K��2�I�O?��Wd ѥ�n2������(uTb��G�b[�$�pyzχ4`�(�r/JS؇՞j�D����0S��_��"�զ97drjP�4���I�~�.9�CФ� J���n�O��Nv�'��*a%xr�CXFVQ�&%�#��lT�~�=y��2h����u��B�
� G6X�	Dס��p\�Z���I��>����,�/�u�K?�(ƽ��P�:m�񑂍�t�#q�"��[-����9�PCwr
�0K���[�i��<��<3.��rPΜ;-�ܪ�4�\�uZ|x��[�Z!GZZ80��DL}�����r�=w�Vؕ��3���N�8��V�3g�G�� ��(VY?��;P3H�q2�=F s!j�@��e��^3�R��9c�,MJ<�j�QI*#���vDߨ�&]u�����n��z=��lQ�wW�� ����T�Z��E�E�n���~��t�߲ۗծ>u�sR�sN��H�A�����ա�נ{�'g���m�Izd��8t���I�gX�]���*p_����F)O���d=zO��)m���{$_��"�;n��>���VY��,��k�14��꿷�<��
9��"]JN�Ҝ�+zx�=�2�k�lٶ[�T���k���2 �e$S�i��X�c6�
�q��R���Y^D�=1>e�V�"��0��ӧѶ���?a�ģ`�L��g"�L*NC�mx%8&�j	XGeY�%N7��0M���*\K�͈Q\�@5����\��KY/��[�}����x���Yv�J����㓲[��/� �g��_^�{D��N������o�EB���<х��?љѥ�d��)9t�9��������[r��Wh���//>�K��n�9RҬ4�q~Wr+�W�
�8�կ�~�<����2?#���|�R-��Gk���r��2���{Ǚ��If(�D��ik��,��H��@���]�'�xB�
�����tOVF'��5���zAƶ�˩Sgd����:Iit��@�ܮk՗�z6��%��w�������X|P��=� e]�G6���u~��(K�)�ݷg�ܴ[��F����;q��<�Գr��i:�s��I��O<,Q�Ϡ�ϳV�tF�t�ğCy������mMx.�K
��C~^��R��KAH�[�P �ˋ�pur	����E��?�_V��OV��屿���2�L蚭�o�܊�Ow��+Ei*8ۢg�K�KRV5�س{�ԺK�G�Ȩh"A����S ػ�0=�DEa�kϜ;KQL�5��g-�� 

��#�����컑_�����&���e�۳���Έ����?+[~=Y��:<9)فa���k@��=� �̙3�,�����{'NG���vZ�Ѯ[\a�W&�![�m�~}����6b�U볲��N�lK�o@�]u�- ӳ>���̹�����.0_ ��	��/�:�_~�/%��5�U_���"�~jBmY&���q��s�(iB�B-��Q�6jdB�d��np��zV5�tkI�L�!E�}R�ם��%Ɗo��_Vg��Q�*ѿ#L�&8g �ޅ�LHR�b"jz����P�~�m��) �� +[�T;e���.� ��0�K�^�MKpמ��ß��}�sq�}���	��ҩN�ڳ:B����tL#=���Ѯ�tPKU�	$���!k��+�:꠲J�fݺU"���%���hR#I�TV��ѲI�]�ތ���'��ۊ2+@�z ^���������
s1R�z(R{X���%֛��k{߬k��V��#��[�l�~;��^��?�4��!�3)���0�+R�$ӂ���]2��#�y0��Z`"|jl���l��V�E���'�I~Y��VP1mҔ���LR��t��l�s��z��K�RhH��CP+u�v훆
ŻB}�FjH���l�ƁFyY�+0�P��iרK#ڇ�KV�9H��g�Sp&-)n�t�D�V���cvD�n��N\W���;�ev�m��ɹ�w�X�L|�gEr�/�B[���{ ��v���sY=��-� �^�6#K+k�P( �я�az��������~��,��'����c'��o�=7�g��ҕi=�YXZ��	��gg�5
�B����Q���DG���c+:���<k��Y���%yK�ҵ����<?�,��KWձOI���g�[z�ʮtȤ\3�pψ���r�\9wBV�V�Q^���<�;u�Y��- P��.-�rmQNj��غs�.[/_��k,��1;s��?$�ߦ��؉S28<A'���c��(g��9f�u�e�� �7�U���(��z��&�O���;����A��x�T��,um`�����ڴ�]����{�1Q�/h�@�&%�a��	tA��x%���?� ���t�:V=�z����?�Ʒȼ~�Y]/*�B^_mڔc
�����g�3Hi2�Л_�ߛ�&+��A2��\�=RW{��@�6ޕr�Dy�Ǣ��<wF�_:O��� {�`�\���5}.K�O�
� ����ZR8_M�%�Д�/\ðS!w's�ۊ��z�v���)�i��Ϻ~�
�Y��>� d�\q�gr�gΟӽ3+��GY��l7ՠ�I�X;s�����T:M%�v���Y}���e��U��WN�?ϳBxE}*�v�z �AW�yv9tGr4��3� �ШE�P��%Z��?�=��n(PQ�*�� ��c��8*w�q�ܽU8R�	��U0/gm�G.]��n�`�/�.oՙ�mL2���S�ME�$2t�@����YS�u��0N�I�g�.��Ӎ� *�4�eZj�X!K��Cɣ�>BBr��֨Y��a�
E��2µ�t{ZӲ) i����χ5����ȥ?�,K�qJ�`���,E��6&`�Ք�~��*o1�W?�kt�O]~�R�c�d�c^Mԏ�Pc���� �d��n�����0�Xt�6ɦ5:�eSw�0�0����� a	BV����s�~��hDӵՐ�� B@�R`ʩ��6�l���Cd��~R�Z�����8H&]N2j͓��d�c�����12.�jQ#���W�S��ﱝ3%1u0)���FƤ�L����GA�4�TM�=Hĕ[:����h��Z��O���0.�aliD	��c�Vu8{�F�.�Eu�'�Ǯ4L\v-Ќ��vws��=�C��t��qS��Cb@�s��$[���n�o��h�Z.u��r_h������tY+�oE�����@.��+� xI��)�M����U}�/��ZI�
dΫs^�@���:ߕ���8{����a�vɀ�Q�q/�#%H��Ok�����<�a\��F�
|z���gM	c��jt���G5¼��׵r]
���ӡ ��Q�g^:*�^�"k�u���lZ#�2����Ԫ���K��xMNS�ʺ�$c|&PKV �R(H�Z��;��^O��Z��J���&�fi-.�Y:A�j]�=�]��U�~Z#��p��g�|x�b$�Ncai��[h�=q�F�W餡��lF�e%m �F�6e����i�\RǨS����v��S���u�hOE9�o�}�����M�O�_Ӡ	X���mI����uO�g�GV�3v��9��Ƈel�W���
�LX)	������=� ġI߲�!PQ(+x�[&�d���&ǥ�w(Nl�Kuå3\��/-6�w��j �]R�U/69�q�Ƭ���SF��KF4�TP�!�>Β7���5��*�� :��1��51����,�������5�5�!�\E��dv7����$}��]���J��U@����l�A��������������C�N?&cS�B/$��`��t��:1 �.��� ¦P�B���ı7�߄Q�"�'�$��C��;j�ѭ*��W�kF�7������o�h5b�����=�e�	���j��Էr^
Q�>�F���K1�´�)ڔڲ��'���c�8?c�]�oݵ�F���c������^��n�8�k8��ĉ0���Ԩ�Zq �U���>��?���r*��`X���t�q>{��D�v��~��D�>���u�ؤ����Py2�c$<�h�c�<UD0:�Gf��n2\#�$�= 7�!ߛ�2j��HF䞰ĀZ~�:��d��]ԩ@g
�ޡ	A�7�H���ǆ�ڂ+�9b�'T�����D�׃۪A�!� "+]��vWed�M6F���z�&341Y^WC��c@^G��ߧ�!�K�K�c����Ľ�
ԒP'�5�)��mFM"��)��j�*7tO�$��1��(J�+Lo^�/r��Q��
�P��8�`-W8Dg�}ff��`�]�\�s4i����sļu�  C�$޺Fk}��'��� r �ӽ���
}� tU����L��'�.s�vup�C���d�{��&ɶU�|��+Y�^�����;}ZN �-�d�-臁c�����vH~}��aHg���cfaQ����0�*ȫ1�2�(�>ɒ&����{Xb��Rզ�Cd��F��=ItS\���uɣ��k��{mv���rjl�Ʉ�� bu�g��뾶^dgȺ�$Si�R�]Y��k/��m\��8��C  N�/�St���D
pO��I���� ;����_�0_R `�dú���+�yQ �KM*��tF+����X�-���'d1WT�s��6�v�R>/3�˒TP��dԡ�$_^�=�N8n�YP* �� $��(����"X�:����{��}�iFL-(�l�dw�3���XQ�.gn^���CN\�L��"z}s��(V)���F��������B�-���㲪6�F��V⬣��K�Z��&F='c�$pV98�Iȯ6¢E޴~�%Ś�.��n����µ(�SfC���̪=�6��R����$�4�
�UW��>�/(S"���v^�� �Wy]�A�������K�+�@
���I)��*2-�����A��ks����^������|�Xar�� =	7��O��#��qI������ٕ%J^���ܷ�K��)� ���,G��������� au��H��3�����&��F��
����_���.��]�x�+�5j��V�ܐ�F�)���fB^2�����#�Q��X���V|�<����믿�6h�PJ_��/ˑ#G��A����������"|�%KŊM�t� hi��]�h�M�� �e @p��-�jb�}�����#/����"E�N��J>(���G��C(2�'�jH�SSy�����bT�L��&e �e<E����F%��ԥH�m���b����ON���9r7#���~^�!G j���loc�)�\���!��}G<�͘�c�Z�6ڴ=�)B�B0���`Ú���}k&o��W�����5�곁�<�Bu�x�M3���y�S1�8ʆ>���Q�Y$��Od�eR��F�-ϲqp��!3���QxC��F=����|Z���;%�]Ýl�)e�c��+���Sw%\�5�ctlg��ضm{�N�۶m�ض;�q�I�6����y����j�X��E��j΋�VZ�*��ʐ�2r�\��j�0��~�#u�Tx��+¢�&��ETB1��Qh��.ag�~H��ڳ��eh�&��J�����茅f�!�=����M���D/����@�ZB%���'���R<��i��$/-��n�G�<�	��'թ�3N����qzYV�v�c�R����"����u���y��|���#��8��"���H�M���8�.�CP���-ιtjQS��i`����5�������@�8�f�W�dH�E.솼&`�%Z4��-�o��|��xС_�Y���1�?$���%)�_9��=�$~t����BC� U�i�wx�i� I�S�p����P������v"Mk�Ft�EϡZ�����/ۉPr�W�#�I��e��9�M�HFc�2~$B1���+>A+{ȍ���hj7��.�Ll~����8�9�I�_����0��ԫ.`�wp=����D����&aE��oC֯rX��ߏ�X���1Xr],P���v�����`V@Y3�i��5�U0�|��DM�u�)ݏ�1��O�� KpH��1R���Ȟ�/Pk��|��R��*
*`�Y;�90=�nƿ��l�aQ���u�[�߳z��;��j�l�ht�FV,�t�BcP:�@جN܍���}�#�~kQG�$Fa�����ث������v�_&C1d��^c�[Fx`Z@ݙ��]y� �B��D���7�]�����B%��i�N	���}נ�0	_|I�,D�}�1mX򲤴��[�7w� �m^��q��o��S�g�������uI�	_?��W���?���M �Ԡc钋��&�ؓ�i�\��&�'�&�S�J��nt�c��R-�c)S�i�aJu"]!6���-�z����De�p�UF������[v�Wwm�X�ߏ�!Y.-S�xE�����UT[W�3�}Wz��~�(WtO��ل^�l��sY��5a���_�UdE9��#t����ѹ�4ٜ�λl�����-w�A������� ����>wb�^�i�^�t�6�vb>��C2�L�-��p{P)����#w�����G��g�
�Uc����!�]�ĕ����	:�X�!��p�&.��[}�tF��\�X<H�Կ��h�$�J->*y>����e�S'��5���B�AI?g����:�*���)����el���7bLʏ�)P0��w��NΩh�f׶R��8��T�����[U�T��ʱY{@��U��D"�zz���(}s�5�>��LL��%;�P� G�ٿ!�~=|t=|�.���Asٷ!�1j5cxe��Y�O�P��wэKqE�r�E�
�����('�Ч���KH���pTwb���2j�,�\�a43���q�T-�o���fXn�������<��0��0��P�t��-���J[��Z`Y�O1Y���ڢ��hY���ǝql1����p\�Z���33ֆG��zhT�p����J �i4Ne�*��!�&^?���slIN�@7��A�`�oǡ���Y�=�)7�qk��cK�������*gKmm�;n��,��.�J��L�5攆��:�Y�A��ş��� �T}���H�|��х8���	%t6��X%�e&'Ӣt�V��;QLޚѳT%�&놚F6�ꭘ���y�0��1���,�m�S���-�\��@2E��L��@:	��i�g�*��yȐr�Ǭ!J�ccٺ������խvJ�����@v��04N"KT��X������v �����!� �����_��><�B#��@a$8
4�	�av������M�d$6�uҨԆ�T���[���l6�*h��d��8pEJ�R��H9���� �]sD�V[�
�`�F��벗��+_�O�mW�zZ3�_������eR����<������������Cy5�6�BHE���V	�C�N�8/C��n�P�Տ2�m,���no��7ez�S��j�~ލ4嗟�
	�,Ci��ss�X��;C��,4���� �+���a*�rꨡ��[��5���%і�u������J�eY
_���2�,�y9o�Ϧ���+��j�ug�����Nv_���b�w��;ާ�z��o�=��K`��$���,��~�L��`t�8bn�6S�/����	���_*KL�v����E���j�Z4���T�߁Cφ�@��^������p�Y��M��<w[��r8je���f�uZsΨ���C�+q�㷎F�K?L����(TG�&B��չ�=�f��D�4�~d* �o��^#磊�a��"������N^L^�F�SE�]�6b:a/˺ͩ�ƨ�d����.�;�*��w�;K��].!�r���0XU=p���Eb��lS����Ӧ�lL�-��^zc�c)Ҥ,��[�� �ɡ�b��3��'��Jx�IR�P�Q��i�23���I�������u�J���s��0g�g`�����m�#n�u!�T�UA�f2���ʠ�}��PZo���������x�xvn>�G�{(�z�b	c�s�ʤ$�><�V�h��SaQ��9�״�Z� 7�do��va3?����r3�C�
�K��O笾��VY�?��CD�mg �q-���So���,�RI�:ӻ�W��8��7�i
�zr�!5��ƿ��� v�7iG�؃����l_�Z�\H������¯7MFVD�K0������+?��(���ͬp��ɚѐ!U�1���L�)���hS~��ߴ��N������l	����p8*+���� �}
zk9�&=�����9G٫�����%������v~1Pʍ����Ja�ezy8�E�0$�5k�tX��5�]��=^��E ;��rM������VQ�f�q�`��9r�hu+�<;<��d�~�HzUx�:���v�zC�V)S��f�P<r����!>����|�tu���������/�0g�~���(l�o�v���g�%�X	��8F`�&z�w�jA����?��y�|#�3��������P��D�,?E#�!QU_��eB`Y�X/1�j҃��^U���L��(Y�9�H�AY���e"����X��0��40��/�ڔ�܌��]}�ą�e��Ln)-���|5�?�n���[��fv)�S�v����Lpeg��%:��B�*��p�8��V�)](�r
����c�F-q�Yt<�h���{�.n�=��>�;�/1 p�+���Vc�=ƅ�vV̄�3Q�!�M���Bk1�@��Jn��"���O?8.c�83�����j�w�M���p0���'~��}s d�G"�t��H��r�W�f�KZ){H}/G$F8�;Т�n���:/m~|������y�h�@���r,�����]�,�X-R�?'��=$��z���T��
�诞=�Vd�1��뉕p%���]k��M#����cj2�����d���-�,���/�I��c�ޘ��	�EX�W)Tʭ<愈c����*�Z��D��WJjR��@T�@?�@!��ϻ�D��{>��z�#ÆHD��^9pz�@�Y)�d���%W�%��i�(YJ��&ǌJZPxU���&|��8�]�i]FE#����Jj���ۈ��<���z������q�iI�{� ����"'��t��텯r��/v=u��'�4O����=s��-�$�Z�|b΢��|�tQ�D�V���'��H� 0���c�6moJ4^�, ���( 7T�P�D��/��Pľg��� �I�8�ٗ^{�q�𿳡���!tŶ�=�4$���8��P����,4��?NS���GK��
��W �1ަd��G\�Y,��a�Ұ\�E�:v�]	{�'�I�f[���gn!��2�N
d�Xrj��ړ��ac��)Dv;���$����"��ڌ5���'^�ϠR��f��K�H�8�����Q�^�2�~��[�}ߜ�U7Q@(GA<g������bN#L�OxIFw�x�4�=�b�y!�9�3��{tSv5.��1������Y��9dQ�ɾt�?�S�!�<�s�U��e}��{�	gM
p�1�l�0�LR�ÑR�ۘ���Z������݂�[_�v59J��Y����KU�q����7�N��X���m���QJ�wl!&����&U��}k؍n���A"'gI��P�M���EA����?�j
���-��P)bW\N'���<Bٖ����k�]`��VF��j���a
9Ji�xz�P��nI���p��]�e����C��$9�UK�ZBS�U��f2_"�p#Vɺ|w�|z�M\�c^DW��2-���*� �XF��Z@����F,'��;���)�e�������0���Yd�n�Ŗ1d��{ʖ�"��!+k���� �b�qS�4�5�`d	}�(7s�,-usw(ʙ
�ÿ^�_�iGM4�O�ω/_gg �9��4��Ojِ��J�vgP"��b�:Q�TmB�����D7�ɼ;�yO0�])��b솗�d��6TN+Y�^���t��`Ա�8P<Me�s�wJ7|L��R�$�g5��Y򛃎�^
�r����-��%=bZ0�Gt����'���I����(�w�ǘ���}�ֶ$٩J��c88ҙl�
�"�6e$^"�alV5�:�������+��!&B�t%��Љ�P��q�-c���s����껓�k��Yw��k$��*���A[6�f�d�����Ͻ]�/W>�\!y��$���1���WTX��ᜬ;���i>vƙ�[�~��/)�<�~����w*Ql��ڴy����9��PpS$��V��o����ג|��cN��G3t��$�.���d-��N�2�;�{g9g5��+3�����*�4��w�X��8�6���.�ۧ[d��V	�z������߳�����*�>"_ƍ�Fk��yeyb��]��T���(-%0);�tٹ*�q�6���g���6"qv�;MAE�Y²�2�8���L����,��ϕ�v��|��@o���8b�(AO��"U;��������U-�]�,��=k�N{���ҁ��n��w�|��zk��S�)#����f�<E��r��h���5��p�	��$h���	��>v�q���mh8��l�h���n�*���v���UR�o���"��\fo�H�ݷn���O��<#E�f�b�9�`�_����	hnBX��cgyz�Щ�-39.r������?+Bd�;����l�� n���bv� �-J�TL�{BL|���[�憯\h~^�0f��+(�c�iKH��z��*h���dk����(#yh�
���zE~�Yv*��aN��TƂ>"4 �Tfo�pݼ��?���X��7C��-B�����~@BLB,N����<�M�Q��ჼHx:����1�{���[�
9����Fno[���栙<�X�Òs$~aB�1�Q1҆RG:����L�,uTA����8�b��v���U��a%��&�QGiI���e�n��� {�[�Zⶾ�6K�zQ�3QN���9�1����Q��\���7�B����#�z�����#�$��}�R�S��18Ň��h�� ����+�*Mq�J4��:.c. ��F�RTɟ2����%�T����7]v�c_�����쓕��U:?�覸�tC�U)��XL�Vم��m �M�ao%���$�.)A������(����Q�l���*,�1M��R�x�C�DҸ'�@���7/�m�����&S��>?�����������+�~�~�U&�dJ�vϊ ]��l-��ʙ��L`��h�E粕�)D�|Yԏ~��%*܏��c��6��$rn���9��>��'/a����{��4�;:|�qB���Z��70�����&����̐�%Ǝwx�z�F�	���N�qy\���ɉlJ�{w��%bb6TgαQ�|���y_�}9D��r�ņ޽�Ìo���JԔ@<�n�������.��H��
a�*�%!�^<0�.����$
�F�3Ԍp;�٧C��;;�����%��nV��iw-
�an��"[����v�i��A�rV��U��ag��$��������h�69�D�$�쏮�f$�W�UvoV���cc���Y�I�7%���9�v���	������ #$�s�:QXh��md�6�M�/q�L>���3B�����7
��RFžDT<���s�N�O:oU�7Vb���cl�`*lJj�{��������c�[��agZr���8�Ӑ�K0�����Ǡ�u6C+M%I�R�������#���C��A�����3:�.� ��=���U�*�
���?�m��DnTw��i�W�E��&�1 �����6���{9��-5

�N�O����:A�"����p#�Mn�[ù��������?��#P/����j��EN�@������p�6�������4?�wT��M3�5Y�����.��p]�����I���úT�d��UEzɏ�hE!`��{��n��Ф���z�z����s꟮w�}���Y�����/���n�尚�u�g���r
2��$FC	�B���;(�������0E|L�R�����d��Z�-���¼�G��}����`�|c~E�3~9���pڰ�|}ɘix�5``CCvxn&P�I☹���lwǓ���޲#�� *s���<�zO V?4$�j�	��Fg˽�g�Y���Syu
�@��Fޙf�S��o�
'~ם=�qn��y�X����Դ����9���iB���&'���"��n��}ֻ	���A!�����#zl�XO��c���4�'�xӶ@�T���w穒�=:ʰV"���e
~�Rm��kf�
!P��%�fo�	�]�+�{ I�?U�Ǣ� ��G��qfv��K�)=�Ĵz�˷�P	�,�$bҭ��H�"�,�GL�f9%���x{q� �e����K�,sZւ[o��E�����W>~���}�����5;���"�|��4�/j��G��4�����z���}���@x�	Ad­?�� ��D�{�G*��qͧ��і������Ϯ�Y�O���P�m�O�#4�,�$5��F՚��B��V�6�j��z(�uM�V�0;�	&S��PR!�*&-�gB�\uݡ�%P�EE}vyMq%!�YU�~��� (?؆�Mt(��2%��j�X�Y�.Z���8{�#X	7/9���[�7R�ڱv��tR�tW Ѱ/�-�>gU�������^Jt��>�+>TH���0�խV��@m�}0;��$[���P�ɘ���-y��l�A�����u��A���zp��U�y�i=ƹAQkt{�%�pȫ?׌�.��)��bE���x!�?�üʂ����Tx.k+)fC��y�SųԐZ�ǚ�k�4(=�1�P�ϱk�l�#��۪�[4��{���ԇ�"�>`��ȀL06��0Fi-*v��O��;h���o�@�Sy���P�O�p�i�
p��'���i\�]��ׂ�'�3⿔�hL(���\oc�{çMs��gϡ��W�Wp�F�G<s�<���*�0���R�LR�T�J�L�Vqg��/8�}��g:�qgN�*�֯ԅ��PH����
f7=��/;I�~�=�� �O�ݕ�&6��-6���ƀ Rgm���B6C�W��.}Y��+�1���.	��<���c1H���+��z����?_��T�M:����3� �n=�j�}���M����� �ǂF���m������)��1��O�*�
"���t�z�i�%�{�ӍK������'��mz%#QG�w��uY���0���E��t_����R��q%٠		�3(��A[���ȍ>Dw�R�0
�,\n� ��BD�:��uߩ��y�p���V�����H�(9�r��@���?�2�#�~�T��V����Jk�p: G^�(���zBvKk����:��J�����Ē�J�T�Ah--C���j�J�'�B����yK�-�Sק����R.Lg��^�9�m�+�H*�N��S��8�g�Mn��ڄ�t�d5�G��mb{(�z;��Xt����ڙ�N�+��ȚC��V�(j�D�'�7��'U��6k�=o��[�x�O�ȼ@>!^�Q< ��(uJO9?�[��Ǚ��y�H 5�W�H� [U<'���]��o���Qb"-;
Zoq��$;8���BSo�Z�,;����n�F��#Wpm��b^K:썓���w�f�z�j�{F�Z �Y�Z�u�������2y\<H1�,�c�������+T ����2{�����q�%A�2�kU�X��H��KPڦ��1�1Q�5�cg�})�݁�N��5��[�� ��5!uBݶj�����2nZ���]��xz�穭=}
"h�v�t'e�|K�Uѵ��KϢ䭨-/�	T�(�銉V#��x��%h���}�DI�w�-C�����c�7�!�rN����Ʃ*�)�s_�K�P��5�'q&C�3�{`���ut�'�f�=�v&_�c��Y�|�gb�Rld��Q��i������Fh��{%lI������J��"��)���0��*�,���8�]7n�]��S�ߍw�}f�x���7$�����q[��GƗ������9w��뻺��%��zT6j��|.w��E�"��ߐ�X'�3�����pHq� �\�7y�ծ�.S��|<���Op�$�!1�"^���d��Ͻ�6
�kJ�?#����![����B����Ϸ}�&�B���N��%Z�l�>W��6��jzwvu\eː�_�W*�0�'Yn0�CGEO%#,�3-;&F���}���J�3M�Oa'qu�^]MmJg�X���oB�m6؞�[@@�K�X��yߊ�����g�j�f�,������0��v;?b�1e�c�C�QS��N0�x�8��z̔]���K�.ª��]~�=�h�g4�/�>�fi��H�����*R��W��R^���M�����Dp���M�=�!YIg���򛗀�3�|��|>�3�O���!/�A��PO�S��p�O�̦�j���G�$D��yg&�v���<�o_%�c3��Is9v�!ٚ���NJ{�2"���y5��!n7�������-�Y�ሖҋ�ZeN�f����z&t
�?$��˶Lr���k�~l��&�E�"�0��ʁ�[��3~�Rq�m�؞{�L옒Gb�f�
l4}���G��s�n����5�#�:+ (�HWu���
�e?�saԶ��"a����9�VLGcYgB�J�?O�j�L�V�OoK���M����t^:)���d�K1���ZQ"�{�ゅZ9���bJ?'d5s0���E�%L��G��
�]�)-5�uF8ңr�`:��L�����O��ݟ��2+Q0�	YgOK� ��d!*k��3��8L>�r�W�/���ȋ2Ge�G��^�h@uE�k�~OZ�b}�H��L�Y�Q$��ܛ�iqw��e\[2(�[�\�����6D�Z8d;cY��BߔbZ���c+]Aي�G7=� $�:г���,��uim�#[~hjlP\:�D!�21	t��� �֓L�'��F�՜xU�2[-����� �c{�R�K�c��x���5ʈ~DcU�0#"i��VA�SW_~��D�=w��
�A����!Ǿ�(�%�ψ4���5�K;+�(g����H��%��3�S�ᶏ�7f�'M�$��>�t>���4�YnG/��i���~���
�we���Z�E)�����Gy���S/�AʋV�)�y![*EAv�G��LU�}�7([�>B��D��CV�ҿ��~�IQ�U<�l����<�\��/9'��E���#�F>fbr~8�
�j���4��̆�UU|0(%���A
Y ��P����*�oJ�)�l������rE��X�j˅����)��p %t_�u�_�~��KX����$�ęC��DB������S<��� ޖ����) ��ҏ4]�R����g�j=(������r�mv�i;�wX�Ȣ�t��%��{�7���l��?�;�I}Gp����J��#��[xWl:X������s�`�&x�f%�Z32xxR`��'�MP1b��Ak+їA;���1�*�l�w59�Ml�p�t(-�y#��2?��)ݠ�i$��6���̅ǑԾ)Z�pD����1�}�����'���P�0���q|P,��9�l,ڴ���l\(���c�1O��ۚ�A����9^t��~����Lԑ� i��.�MLȐ�
ukaHi,dj2%o@@|�u��^aZ���i����`�Z��%cO�f7�&�� {�`��za=�u�(�N��ѷh�з`N`��e��5�ș���k����X©��-'�R��)8"���;��(�#���8�:v�Uj+�������/�0���-K�W�}$[6
�>^�N�]�7|��m���L �^��6�.�����"T����?2����FgQ�Y���$N1y`Oor�&�KpM֛nX��n�f|�~�,0Y���J��Ć�%v���>[KV@�T�lBg�U�@����它e
�x��p�v�Q����� �iikD�"��f;�d�� 6�`D�g�̃�]w� e@��(Kx�)]��ܕi�P���
E��*/+��}3��ݑ�vWW��xvd	;N���i!c���P��B�&TK�)KT#i���Q,��k�sX[k6���N���&	t��WLA�G
7"&s<�h|��l!�����Q��Z3or$8�jr6�u�������-�[��;��f{����k�~ڦ	+CaLf*]�^m|&9O993$on�VU1�h,�ٝx�	����5V]����������E�u�a��^|��LO���(Zk�}�EU��s�q_��1�2'Y�*�r�ףw�d�a�O}�D��iM!vt�?�g�F��Ic�m����CA����4���d�
}ǿ֥����F뾇ͻ�:��,��A �S�\]�!'��b�����Ǽt�y4�����[�fb�{iƚ�XY�j���M���%� _�'mG���U�����Ć��H�ܽ1��$0�Ӳ�vMt��6�H�䷗ܽک�pQƕzC�\�<��X=�0H��(��<>��)����n��Г�0�`�Q�4Ӱ�<�YkwBBBG�-�#5�x�xjk.v6_��bB�Z�V�Fw^G�*�֑y�����Ҵ���hT�[��<T��=?>�$z�V���aƉ��ӟ�x��iǍ�*�J�K�3(;��[
\��V�)���ޘ���~A�t�K�֭��?�9���V=�<���>�}~Jyӱ:GQ�5�Sox�� ���`��� sZ�J����1e�dMh�>&��x�0P�����������(TA��ldTF�=��Ƹ2�@Nf�j��¹����.ud����!f�O��I�ܩ���0p}JF�*
*�"��:��k>��8"搐�(�V�M���ƣ�W�"(M�)�"le�18�>��0�����i�!,t)��7�V[!�3��) gcj��2Ɓ�U�Vf�~K(șa)��I�g?�DL/Up�7�W�,�0��vf�6�/}2׹h�&ӽ�^���4�p��Rm ���3�B��(��b�*VD"�_Xnt&�՟�x�N������y�҆�O� �X��PgׂNf�a^��ĭV��h��Trv�Xe�)���dY���
���/��E��km4���X�� ���(+�8�o�+&ᨠ(k�{�
a�|���m��Z,�b��w�;�&�΢P����8[���FK�ə��sZ��	A����;��F��e�#4�ްh`E�"��:��<�f#@y:\��¾lj8/���B�HF�Y��1��x�IH��v��o����bӪň�u;ICs��eu�Z�jxV������t#�ݥ�,����>�r5e�na�b��׌��~L���'�O�JY�3��][]�3�c��Ǫ��e�������A��)8��c4d4��gpvF0�Z�S�Cb��])BEr(�CP�ɪR��"�;��I�<r5#�o#����[�T������P*���Y�5С�0����IA�1%�X�"g1�w3��koɈ �~��+�iE��?�!u����#I�JE��^	x64��=�4���w�TZ���^�oh�ZtOV�`e��C����.��"�|�q%��$g�雠rS�@�ю_~�Y�{����e���7ǽxF�_ଫ+�JÖ%�#����J;qo��S(P ���5!{���5���}#��X���.4V���(����h�u��L��g��.,�#2�?�-$��9q��I��>��J7�&�|ڕ���Z�)R��g�W�taCv7Mv��1�� X��Kw7�0�����WQYG�u��
n�w�薨��9�%�TW�<����?S&�}�����R��ק��-���x֎}�F]}��-��|ȝ�g+N��nu��_�����1���Z�q���kpq2��-����E�sŦ�ki"֓ �]�;o�M�x7 m!�MЭ��7�D� ��7��M�85�$����E(οM���A���t,I���i�I�/�d��� �<�c$c�oYA;C�8����!Z�A�e��v"�ޣoH�֜�$����d�c?�饹��'��۶��.'��� �ի�*��upF�l�12���~��3�"��'�xѽ�?��w���ڎ��2a���_�o�}����]q���%п��]p�M|8oxY�i�s+�i�1�ܕ��������g������P����3k�\��fC���B�T�s��V�W��O�Ԇ�0ٚ�6~u�����I�4��M��,�N˿�V����	/b����Ă9z����*h�e���C��U�˶�Q�tP�d�%�9'���ZسfB����d�bIp]0�P�˗\@.�<o$�!飘�$K�uF!F��č��I�i�bq� 7�+�)�|�����?0������0�%���*��`6G�:�y�Z�a�o�i�_��0f`�N�G�ׂJ�QO� �$�K�IK���u4�Y��dO�2K��8� 
�s��ͪؐ��
D��"!U�Ce�������U�=�.�/�v�~����~�����,u	�s{s��#w���ν���y���1~�%�e�cb6�����M?�/�W����6r3Rvw�hup��#Ű�}/7L�4JL
�m�^�����A�_�s:d�ւ�!���M�#������B�g�(��}3V�������N),�C�v��CЃ��M��t�Q@�&T��$���c������4�=����/���������r�T��}�ϫ���<tYj#k�/�^a�-Tk�_ǵ�_(?IyV'�~y�V�YI%�z1���PK   ���X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ���X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   ���X�'k�  �  /   images/e8452abc-1b33-4025-a556-b46ce3c60df1.png��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[	�U��j{���zI��t0i�D���H$��3g<zt	G��AFe���(*3"�":.�
!,*[�$d![�ٺ�I��o����ߪ��@:�%��Mn���������zo��{r:�P$�����Jv�W��!�6Uuį��뚃�I�Op~�/���$�v�a�Pw��6�>j/��n���G�6�Tt��}l�St��~�S�J8���'����ċcÊ��h:��<���c�$�	�4@��}WM-M;0��Ј(��n�D�:��朵$��x���D����!G��t?���k�~�����]r��4�4��5��&E�NxO��i��}��\<�a&�9B�o�؈Ӹ�>�3+��ry�]T���C�ُ�ˏ@J�ìkA�e��(�϶��Έhϵ��3!��ܹ�!U�Ba�]�p!M�͜�'�Po!�8�I��sm���}瘊K��de��`?Sk�����^����i��P�"���b���LD�	��0/��ٔ��LB��:~b��*4��t����9�ae��"�K)Lȸ��t�y�GE[�e�I�Nc�W~d�⿎L}�B䉯���\a�d��V���5lL��1P]8
&]h$~�]�,��D���Wqd���t�p����1��jS�_[!b�tϣ X��B���cR�Z`�<X����2Ix��<ԧ,B�$1g�x��qV�.^��H������'N��B>�X�Dm}Y�ܰ�w�G�'f�y��h�2�r9H�	��gM��[�K_�aȧ��R�	է�fT(H��4 �^�&��P�j(Z
REx6TG�9LL1�z�RqZz4��A��"���jנ�	�W��U.P��m�ϩ��% W���ʑC�,&�� ��n#�D�j�Y��r�n����{�}�,`�@�f��I�|#̴i-T3n\>��щ�΀E�i�w$��� fϞ�k�����'.f���2A��A���~F0�'oCJ���(�Ť����j�Ѯ���h�v2�A�tt7��ۢ5I�+��>���� l^�;mC���v
%Ocڇ�N�!=z%�1���DL�����S�v���(�l�EA*�&��{;��ͨ8�MN:1t��P
�;��D� �?C�Waeft�Ǖ4�E��cČx@#f88�ȣ�&���iHU�h?�O?�$�.\H�I��4�2\��p` �H9�~�s;��/����a����0SK�*�a}V�g�F��b����&b�Al���j���A���o���	�]���VPtG�_~Ӆ�k�m���Q��`�ԃ�R��k����ކl�h���|F�5�����=�8O7����G�M����.�@�������G��Ryt&Iw؄h$	��":�%�>�Ïko��h�Q�1��H]y;ꪪn���K�޽�q0��Uo�`�RF����V�H�J�O�IT���Q�OP���$��"�
�L�k)/۵�8��6�I`ŭ�G����q8w��;y�y�������0=��D^��C��/K.,��E���4�T	�����]�<u�.���!��XJ��������7L̲ϙ�2����/���3���Y���1�"�L���%?_؞S&`�'��z�ʛl����9q,�"�d|�T	ӟ��4>��@���z�ۻ�%��!�m�w�Hr��A���+��@:�����A|���&�g����_��IÞ���u�1�y]���e�#PN"!�Q=�?��*b��;���j��i��Sf�R���F���,�aS0l��q��ڎ")(ɒ).��֧���p�Dmď�����t�CUdl>�Ep����i��5k��U��/�sd0��cv}�����m��xlk~E�wT��!̌A;�����R�o�pѠ�|-�WJ�xӨƄ�$:���H��X ym�E�R@��"����k$�:s y����1��fƺ]�8�>&^k�ϒ�G�X+�j���}�\��1�9g�^�eTo�z�`��}fnH������[qo�u���7&p��,_�4!E!�@���-˂��0MS<�w��4���4#&�>g�ْL1��]d35W"G��5̫���v�k*���֭_�K�/G�$���(b�`��T^����ά��C�;C�R�׆��Л"�9�Ag&���B��d�������4MS!Z]�444�
݋��ATWWc�̙hmmEKK��$:::��da|r��Wa�Q(`�h��Z��[�$DolCb������"�Yd�.��PY7�v*++a��0�����Khj�~�k�-|{;��e1C2��!L�

�V�x�Ј#VD0��e�SIn���V���)��kjj�`��Fz��؈T*�={���`�����*��ӧOǆ#q����c�k����y�SEL�H]&�%�m�=C͋������'��ޡ!��ރ��[a�*q�3����%��U����i��r</���l�\�.�ڱ
�)*&�E�ߧɱ:b5��:�Ţ`��g���+W
	:t������/b���طo���3Y\gFB-Y��&���M�@��*�dڞ>pS8�HӸ��B���a�����+?F�#�@	�g��N? 
&���h�˒</�k�M�;�I�ò��Ff!6Oɴ�
�^�7n��ȑ#BE]v�eصkv�܉ٳgU�u�Vq��ö�L[&~%<�� �-%�7�I"��Y��
I��
RY��W![�`���~�0�n���/aْ%�����˪��W���"����'�"�����F����Q�|j���N��Z�C���ǠdNڊ0CX-����Lٿ��f�Ē��mmm�%����=y�5Va����TY *Ո�
�j?yTgTI9�.�>2��:��[!�Ůh9��9�%��S�e-�z3�;<�� ���ݨ�6�*�Y �J���͛�x<���.tww�w�Vx��ѯ������8�3|4�O`*���0� �xW'�ɡfV�D�qp ���]��KR���6m:ló��a��������J�A��]/���"�ߎm c6��1���3��[UU%ο��jkk�!����bH$B���L{Y\�Btb�b�؅̈����	l��p2��$��E��� ��]���[��d%2��E���Q[Uq�/�o.�UV��@-_0����w�<<Sh&�0���l?]ac�c�aJd�ذ�
c;�##W�=X���0q�3���H�H*~��p�]����ds"�ۆV��ae�b [Q:k!�W}�?܃�tF��H_rl9���L���{�xte݄w�F�xU'��J�H�H8n�$�P��]��e�a/�$�y��R�2
KP]��Ϲ��zT$��y����Z�.���B!�-"g��/=$vk������G���éK9!�(/�=OpM�-��:VaO���,I�>	/�\Ċ��w�Q�Q��R��Ҕt���έ�A.o_�("���_{����}��f�~UxY%o?Čס>�?�{�~Z/���q��[��!��ea�Y�k��7L�QJd[.ֻpsh7μy����E��f(}�1¦,$r%�0�"�sk�¸�����J�w���.���_}��H]/k��4��T׌�6��؏.+�K��g����'��#��c���y�`{ ?�R�_T��X$5ў�(�.��l�Ķ�j�^�C[_��T=�����5/\��������tF}Rz��^� ������G���<E���L6V�L�퓧������;}-^'f�j�Ϛ �����EBIlPu�d�He�����8�)�𲊤�T�!�����?q�w ���#b�4�}b?$������p�|Z�P����8ht������K�N�ca���$�r�֏���<�t��,bjysJ<#��k8r�LT�,�h���y�}���Q,oCJ�_>4a{G�n [Qj�;�V�A�{�&�
U#���Zɡ\�����ק�e��gޫ�]C#�a�E���ӝi䟸��xj��` U<=b�;��7��[����f��:-���D�������8���i�i������.���7�v�rkx'��y�	xp�e=7	/��H}��I�v#u���҈؆��_T�lV�8���b/�S��i�dJ�ѕB`�;E|���t�b�e�q|Au�b�w0��f�3T��e$��׬���c΋#�s�nO������%�І^����\�d{!��Mqa�_h��u����"�4U�9�B)ً��F\r�%�'��
��kXa�&0�OQ]Hu�H.�=�c�əʹ�*���O���"����u����1(�%�"ͺ�3!�&�� ��V�~�Ex]i[��i.�[_���ދ�+V`��,�C��s0w��7�r�8O.2QC�	��/k��/�,sl���-�.X��Mq3�
�K�HNID�?�^>8(��_U����3�\9H�D��k��{�݇������-!�`(�_�����.��D�����J*k�)TV�038U���������,�����Nz۽�%�G���f�7�D��؉eq"��� ��N�6g{�,�Y#�!�Oo�}�ń�Kj��a��hy��]E#��}�uw�c�j[���_ �ę�4T�\�=uB�M8>l(5��%�&v�!�:�?�;�fy[Z�3�%�ENw�?�ݬ.80s�|���{~/G�!�a�����
Q��;q����#��A2�<�1Ln��a����,�8�p�p`J&���?��B�``�t]߲C'��v�Z�>D����ؒv�~X/ݏ�?܁���U������xO.�b��)J5ᛄ�§6>(����	o�q|�y�J��~��(8VKK���و�l,F3��S���.��	}��, ,i|�y��y��!�N�sv�z�"�N��&��k���l���a���z��#gaQ�ii� ���K�����6ࠀ�IZ!�#�l?����1��L�$�RQ��qR>>�ʛ#g�X���:1�[��&>�j��Hö�h~
2�e%&�e����P)��u�Øla���1#*�8gh&��
�wh}�P$Q��SDJݫ��d�"$	�f�CM�6(���K(�"�22�
��W@%��I�p#��C��E���-�?(#�Ȟ'ٌ����.t����)��B&<Z��:�'=~��Y��.�U�3�����!�P��yc�/�o/�]�����������I�nTV�q�G>5{�������pw׎HȤ�����>gP.V@|` ��r�	�L�0����2��~K�+R��"hOj5�U<X��dZ��O�L���:n�Bm��d�'��T�{��M铿I1�6[��`sp� f�DB�%��/#N�����a!1n!E��`��ջc=�q�}�����d��\���yMu�&�eq>kX-w2��b̟��HB�I����f��ؓ�ėV�G8R��FVF{�5�{r2"�#v�
�9��mT�H
�̔B��}ҲX�C��I�o��ICn�N8�.#k��;�2>�����6��Ǳ�`�!i˅� �]��f��q�](o��G����9�e��:Ё�S��*��b�|d��E���םX������)�؋)YT.<�<Mܻ�۽�M�W	�I�h�{�X�3��wƻ9#cS�]F|��w*�������������G������ß��go=<��c���79Gu�T�iT?�';T��G���Cf/�jJ�A&�	X������KD��'�o�
2�Iˆ��    IEND�B`�PK   �X�X1��	B6 �8 /   images/e9cc877d-5fca-438f-8a74-200c5bfeb6c1.png�zcs%@�ml۶mM8�m;ۓ�ض�Llg�ؙ��ę8��~8����S�U]ս��U�g���RQ�AF @ C��.�� >�epn�_�&#V?KtF&+�M�����`Ń�ø���Ml6�;�X�{�	V
�lBzOn�_yE�����o��Ϙ�F3�~�%�Ji&=,{H8F�����\�~�޹�kȻs]'DPЌo�$vu�o��|�+��K�+z�	�$1�I�((x*��Tl�ԅ3�.��rT�������!
�?����K^%�U>����+���h�Ԧ�AhX�Y����1�O����ԉ`i��\�=���J�p�փ��\fQ�h�����(��/������"E�|�Q�<�f_��a`a�g�
&��h��ĵX�63.��;�A<�;�|ȒiI��n�+#�X���=o���7�����i� ����û��}&|v⍤�[�GD(jO{�O8�>����aح�f�}�%����#P��+��kz1�f.恾k����nt�5�sPf�����3���Y�쏣ؔdA��K>���=�^��Z�m�W���c�ՙ�쵑�5TK}�|�O��A��M�m����f�!7���@?<���%fA`\䲔�mp�1�WX������/'��Ǜ����~�WG��X�1˼ࣣ��vN4����<(񉡼^��U&to�݉��O�z�ͮ�D㉭���L=�t:�+1Jy�JBW�w*IM��]�������T�̿�H�:��R(�׬	6?�^��޲�f�R�{Z��ZIp��t�ŗ�[Y�W�#��gWX�f���	��$*�ϴ\�߼����/�&@��Y&�s(�t��d_�͊��>���GeK��% �J��Vp3��bH������Γl�%u:�ת��6�>ȥ��s��)�����5vB��6mp��8W���VN�v�wX�g0����>S��C�9�P�Bc��Pn���صVפzl9�o�)c�?����<q�ԇ����),��O�>ȕA�W��po��ò<g�������=��_�۵������+���V�ĳ^@�5@X�ķ�$������Lժِ�yP.�K�qĹsopz�2�E҉o�Tv?��qiQ��@���L����|%@����E|�y�s):�.ʁ��bf}�LnJ��C�����@��+�T@�lK�́Z�����{K�-.���H0�[rV���p\@�%��?)[j�8ba�����5�4���UVy9!�u����Q�(��p3c�m�<���Ҵ,�{���Vl�ǅ���j���~x������lg_�'X�o���
f�5P�[WDy��ҳ\�é�)��Q�v�i����cyx�6�y��[���)$2_�@�k�B9��ē�6&wQ>L�ѓ�"��1Ė��3��}�6�������A�ޅ}�i����W}�E�X-D_�¦4nޅH.�ͺ"��T 	Ѵ0AQ+֟��Bn�P��0=i���x�g�֢�	9�ō:����#���z� ��+��G�	3s�g��{����j!���s+��܋#P����H��f������y�Q�e��0 ��+�lp�[�[?���=�"�;C�L�V��q��.BH��a��Q`�|M ]<�`]��ؐߦ�ل��yb�v���V
Ó��ʯ�B��M��su�Pzh���>H���3��㴆܇yݟ��W�O\������܄��w�g@�3i�J�RR�B���BMz��<&'�<�sa��� �� ۼ��ᛢ%���$j�<[�J�j����sя;��"��8�%nEN�u��D%M^$�|s�lӬT�J�[w���<�b�l� �մd�K�uEo��C�=/[��y�+D���L	� � \5"u����2E3��@b��F��ۓ�n��&6w�d���D��x�is]�S���6��x́y��4[�&��+{l�U�p#���("��*)"ĉ����;�Ͽ�//�-��,��ёʸ��?��dف�&�2�
�>�W�i����n7/4��'�N�;�i}ɨn���$�,7����G^�1D� q	����.)��FY��A���+����`�0e��� x�f��H��N1���@zP��y�JKA����2b��}!��rR�!Ş���h����i�%���"�7+��s3��a������)@
�v��Z�D� w�S`	Y�9[�/?B��:�OG���w{��ox*1Wg�]�o-Щm͝��ȹ�^�������}�r.5�6��q�OEo!5kVz�{ $��u�t�)�r�,����ي��94߂Y^�3�I\���D� �ݷ���ӟ���T�w��
?���� ����ÙyHk�׻l���m�UI�[��
�ϐ������!��QD�"�:w�Œ��ޱ2Ш��ƅ��~"���6M�,�Li���fS<J��k�q���Zf��v�@3���,�<�������#�?ó|�
K�/Y
��]�4h�����s�&��[�-営�װ��9�� ǗG_�Z�sE�%�-.�wP�L=����&�7�4JԾ0��|�Y:�o��@�Tf��#�'� �-Aa�-`%bl�DN�I� ��A�쏚n
��i�V�:���&/�]���ȩ��@��k�Ʈ�,�w���+2��g�@�u�f�)�Y�;��g��4xtl��K�wp����e1��w��P2e�naIED;�w�4F*��5q������~��W�"U�GW�qw��$�)�WG�Y����[v}n}s���L/':ķ�z�;�+�msL�>Z�LL�`&�Qb�0T��X+�{&�����b��{����~��Lƅ|.�a@N�C��!�O�I**<�t�I�W���V*�BR�v\�kn���r�"��ߪ��7�ҙ�E�A��%q�Y���4du�qx�5��p ��C� �d5�#(��]�|�'���ٴl.#��.����	��#�n.�#���:A':H[a��V�H�T\�(l&a�@���>�`���!�� ���#6}�L�2�@�A�n���iGkj^��\��i�vLt=�;�ԽR|���,ߦptA�����A(��e�m"/^(���D-�Υ�%����];K���ڃ2�Ґs#�m�S�ؗ�<�C%�}��#��w�� f`3ݳ��~�`Y\��F����B�6�@�eǲ#`�C��~���s�r�t�kՋ{*s	f v&M�,"&�1�)E\ҋ��:�	�2x�?��Z�q���%(y�$�ĸ���i�;rͥɞ���QB���g�����������[�B
l��Kwt	�1���d�@�;;u=!Z�=����ς	�_d �3(�q�25�{]z�.u�rҎ;br�Q��_Lsv�
!3���Ee]F�/,6v.h���'zu	`��.�s?;N.6&�mї��\N�[>�_,+EU�	�� +��;$��ċa���ȟ��}�3�5�=g=��E�G��=�˛.�Cr4c�.H*�+ck�O���� ?$��^nJ����������0�
�~DC�s@�,=������%O&ɕ�j]��>7���͔�q��2]K�͹ HS�a������3��ͣD�u�SPP�ݕ!8��>X'qntU��S�)t�7l��������!X?�<�t�0�pYƦ�ì����n����ڹ�Ϫ r�=!xah�ӿiɧ�2?f�cbO�s���aU%������ڔ���ϑC����O��H:��p�t9�I3��ߠmj��(V��'�5�7t��9���vG���z��6[n)y�n9K�ن�*,G�FVb��c\(���,h2$���,X��/5T��Xt+����9h����\�(�d���鴣:Z�g3��3Q�IG;�y���x�Y ���F��
2�r�\=?�޸.g���~9�r�-T
'���q�rݘ��� 73�KA�>�?6h�K��W5:+���P�Z��e��I��|"�[�*�A��#�u+l�m�$1�@Q�7 {́���9��Z����,�Y!C�O�*��#��,4�}=�ϭ�^��j����I�d��#E�F��Y)|W��X���K#�vs�q��8<,u���!9��`5��Y��;r%ɖ���}�G 4s�I��$�,H�;�������҂�wR�xm�C���.`ƻt���2��feH�Z����Ӥ$���?�fO'mG"I�#X��4"Iy�l��������`��rq�	�_�I �-G\?�����΀�5%���V�H�(�� se�S����SF�@����Y�M�W��,婺�1��7!���5yGF=�0���V��O7E���9��
�ʖx�6){ٮ�c�G�X:��ܶ���0Q�iu�xm���ͪ���]��됴�2W��ǧ�������;�""0S��6(ik%6�6��M����zru�Y�����x�9W[�.�:�xpv%ZY��"q�t�cX��9�i&���:�����ۿ���??ޚ�Vޜϑˈ��5���hIM��h�O���W�-�F1�}�4����km>ݔd�r�'/�&���=���Z0ڡo���^�l;��%3frZ�F�RZ���HhIn�r#2��4�^X=�9�e�4lP	Z錯ﯧߡ0n1����A��(�1���kWݬ�����(Rv�(^� �r.����o�8���q�	d(]Q�ך�g˙��8;:^�d�Nr��|.<�J0JW�Q1z	��,�u+۰��N��)+j�
�tɕ�w�]��Nܻ!� e�9<��U�����b"�^�qM�\FŦ�]W�$|�fTx�j�D��\��"�BĂO�p��Tpxj����n��}K��x���]���/��.d}��$2@N��T�tטA2p2Q�nt�+<�Q_��=���s?��I�JͿ��f�n��*���/��kˉ8ԥ��d�v��p�ȰY�Z�8N�k�k�T�3$�)u�p�25�g��=ڊq�yi�_ū9��'�&��,0��9/��%I7&� �#"8���Ix��7��g��wKu6nLņ(�V�ţV���5�ע�t?�6uuu-�4������pQHA����f��\1���T}1B'�1�� o�AC���TK�l";��o�m(}u�*� �l�����"c���1Qq�C��[�ޅ��/��c��u�ҨK�al�s����EU���|�	�nZ[�<2�8)�Q�*�4�_̮���a��
�c$��}��灑��_V)����2��l�]��	����f^#C�j<��w��^�z��>� >>��VU�]����X�Eh��]�|��V���������xE5�3�EO_A'��+��h���e�E[[G}�
���*�5�/���h2W��諴5�,cjg
?�m����_�GB/��x�+�V�Y 'ˑ��~|ˢ?�G���B�fp��	I%1��ԟ��<:�(dƐ���ReMl��ظ�Bw�&�ܜc�y���h������hG�)��@4zG<�9d=q�NN�����B�fD��9�4u�N����ou��x~�H?���� B��H��iq�+w�pb��f�#��x�����Ӈ@aaR��F��F��	�.��2-�|�L��F2m�\5�(�2_rW6���|~�e�*�XWz,C�.bd��K[�\���ɽb��DO �iϋ�u�.��{�y9��Ď����i��F�uc�:��d��>>�	Ytܚ�����^�Q�� D=�J�qh�K�kg�j�w��~�@�̙D�z9��\ɳZyx���HʯUݑ��_|�e��UX�(=p���s��lM$n��$��4��@Eu|�X��49��pGөf�=��0�DBO�ƈ*��7�_�1�R��o��l�tO��	�9�em��d�?�*����e�O�m�蒫��i�&�G{H;�)����I��d���ؐ���<�A��>JK��rd�A0�R��q�y�=���jZ'��<aUF�E4����()ŕh9��ɓ:U"&""a�Kt2���K�Tg
VT��d#/��h<k8��Z"̉1�꓃ VG$�Q��XE��0���ƢW)����Z�{�癥�ʀ
[�����~Jj,�M	^��Jx�wEP��B�0� �W���[gg�nٓ@�.�&�v4�y�u�/�m�8u��i|�^�]����9O��u�މ��W�`>��
Br�uO����ٟ/�{�Ǝ�a���M����0URPܯk��K@����jL��$6�Zv1t�Q���!�mZs���.�p)ǒ�IEx:3z�*<�.4�qY�W9H���1F�R=�M��r.l���k��0Oa[�ynD;O�4��p�|\-�PӖ����[�[L �kċu0���r�e�ܭ��r��"c�1XJO>�c��0�����#�L�-�Ҙ#/�g���� �8��"�T�:m�{B�mg�9��#�K[ ^�G��%^=��_`c!~�*>��p�"� �� ֆ��¨��-��<�7�J9���<�����H5[~���.6F�G:T�5P=���G���K���=,)$z�j�P���U��\�C�:�>uNw��+�����c Ś�I�]��m>�O� -��v�]D���:�ѥ�$��,3�!���R�ӡ�,tW0V1��6�
�QW�(�y|n`��Q�OXE=�|6�x��]�F�Y��Dw$'n���P���ڸcc�G��B�cC�OTe�ڌ��i��?�VROS�^���n�C���f�`�S�Odo��(��X�(3J�Z�.�zI�z(�]}�-�	���G�Pa�P�!F�[�4�r�斿1X��̴D�[���m:�� ����Lp��,�Tk6�wM��`�:k��C�${�ǡ4��:��zN.j\�F)-���+ڠ]��LoL|�FF@�_�����@r�Y�Sn	JH��h�i�J�z����n�ͱ���](K4��j����v� �%u�Y�	��>�_V_U��s���P���6$�@����W�F&���Y����1�B�ã�]��!�NH50X��H�S����!8�Zp�?k2��V�up�7�Xz?�w�p�a\�7۰�lޤ_�]�AA�����>�wIư*��s�<�w��������_�?��p�U���/j!p���9p��H��ze�>�\U���{��m�	���@^n�'9�MpT?���	��̨F�C�b�UȮ͉r��N�\���uBqr�E�jM��	n��J�a�������:���L�S�;�@h6u �\fv=�!kR\݅�:��"�.�{����zU,�Ml���d����:���KVu,�?�B������"l-w�����Ͱt���ԁ�P��l��3gte	�N��j�GqZ����M��]V�qj�ڕ�AK$NJ�c0���	3�D��^����ZJ�ﳮ[�\��[�L�%��`���6O���ĩt^����W]��:�CN�l����wN�h��)4%�my?�j_}:�#7��w��dV�T��%B�(�C#=p��7B��H�;7)�{�����#�w���S	X	�D��R7<Bb)�*M�&#{��½�l�Q2�!3U\���U�wN����!=;8�ʒ�q��|�@i0C�Ɂ9ȹ�+�2��u=�?Q$ū�4��E�2Ԯ}#L� 9���S� ��$;���)���5wi����o.����|�Q&�=�E1yd��y,11��|���+o
���@w�N�o�iRRz�q,�0Ybge�F/3?:Xs���t+��l���TB��rr��xJjR?���qM���LC5�ۗ��[Ӗ]���k�jRk���l�2��l��2'���i�����-�,L��cȈ�Zm��QX&�2�l�I[�%�0��z�g/��#���=�{<�y&* ����D1�97�����up_Zr�9g&�$滘�A�ɐf�n�Y:�E�)�e�Z�� >?�Q���ZZ�ڥބ�����	���2bC�������䫂��L[Z[�Z��;'n�p����mQD�@3�Y�{�w/{�����f�uz�+`�i[�|��˕*D������*��*5閊ޢ�qe�
TW�R7ys���͏�z�
!Nm�q}��'�������y��"��U�:j�/H�d�XTƘ�9�)'����]���bK��Ɗvܪ�M��0k��vp�C�o]N,\%eA���Z٢���~�|��Sb���2w�$յ�鶨�Э{����o�Ns����W�0���܍s��׭<i�SH>^^�����F�	��ju�l1�ٲ�{&=���3���	d^l�ـ����nQh�yU:��o���r��%�*òc\���1���b��t�V�UY��#0�����&3�[HUm�p?2e�$�:�i�Ϳ��>)zn��4�Eć���&�O�^j�ۗ+��iK)�O?���G12�L��(��%$t( ����S�Û(�U��ȫtQ���3��w�I�P�8��(.�� �*�]����I��@ǹ��7ܹk��ں���v�C���Ȫ��:�X�go���$�N�V�G����$Nj{2X�	�챠��x�F�V�8��%`�{��4}�{ڌ/����5��AIC��Ũ���ص�·0����Y�ӮS�=M�����%6���.�A���_O�dĨ�&�]DK?IJ,fo/x<�qUo��r�Ĉ�E���b�������,�j���?��9�wF���֣^8�%���������&��P1C�G���'���-����v�-�g�R��[,�u6CN��ڹ�7,���{��U�$r��m̔�N�t����`��MA�������!?͓~�I�������iI��Y�R5�|:��@��u�EB�;����Gˠq�v��,F��Ymc%�?������E��r��"���Fy�����oW�c�Ƒ^~��juk/\���	tT�������P�v�1�L����h��I�@�2��ӂ��l"�����L�2M���3_<�p���?��o��2%$e%YdB��Xf�T��b�qW$z��,B^�����Gf���N��v��X&<��:���V�
�����Pʢ�`�5�]18,�qʊ��{�zXӷ�ƚ`��L��M%C���{͞����s��g���?� 
���^��u4��|KU3�1�0�뤠�q��w����j����Ȋ��񰸸���n,��\�5��,#�V�߰� �y^�+�!II���]���Duj�ӽE�����j���%�d;e]&	K�} �F�k��nn�ߵU��5�>��� |���`_&k��bKծ����>�)���F?)���"n�qqL���0+�|�º4�%d"�K҂� ����nL�R��aR�B����3N�N�ࠩ��o�F���Os�U�\�|Y9��eۂ��� ���r��w9Q@Dڤ,�5Wu	���Z���o�����?S�<��R���sy8��+++�������-/d�8��Q�A�C��@����H
k.������T��C����?�\ԪO[^;q�O�T�Hy���hU]	v$�4ԓ�r�s���:yZ��gg�-�;o�D4���ʴ��r`��D���R5J�r��������u�<@x�g�T#N��]l�L�t�x�����r:x�~B��l];��h�]cp=+1ն�|y��]~���!j\��_".��gf����������<�'Q����n7����_৞��k6K�@�ڙJ
� ���8��A�GG':�j?��$Z�QêP�z�Z��.7K��Yy�8#�{j�vmq8�8�(���2-a�jc��2��j$�ţ���E���_�W;`"�t�qڥ���N�k�+R����� ��{xH�!�j�+F�Ą+��eq��,ȕ��x�pft���:�_ O�j\ν_Ϭق>�ku��ܩ��YS�5�`�-iR��3�<��&�S�`Ц��T��]uC��9m�g�����߅��Z�^��B؂ҩ�F{5��w��[Y_���xw��{,�`���S0�����)����SB��.���V���2o(����֩�Ol+a
�K$�zzВ�wЦV�b�!�3�W�}Dށ��N|��V�̾/�JE^K����ZpX�_X`Q�3��,�y����l]n��2����L|�0�m�� ��T�m���%=G�e�٫c����U6�@��v�o�j���yU�|}}��Ȉn'�����au�l�݈т4�n3R�V��c���Z���Ec������j�*#R��O���:h�ӽMe�Q��銉V3�9�˵����|,T�;�������L�Q����2*���������U7q�L�������<�5�L=t�hxqu560 ��Z��ɍ�l1��t�c� ��j8t]�h9�a�@�Z��q�4ݷ_ox�/�-�.�ł��#���V7��h�Xm�� ������~Y��%�s�� l��M88(�- W�5�|�|mT3����!�n�F1��w����b���D`S������%%x�V����pF6�O�6d�6���F����(��7�-}=}M�8�oHm:�@~���å�s>p����V{6�Y"���m���X) ԣnN@ ���.�(o׻��V9Y0ǃPj�F���Ӣ��G�W�D��5"/�����@U�h�]�S��i���4�����ȶ�a�q����X�W������p�F��:yh��?��k��i�t�n�\|�g����Sm���-�޷�����uw�|��8��Q Md<�+�����i$A��o���Q^�	�����(yF�JòDIy�^��G�]���qf���e�:�{ږٙ�s-�8f�	�]�-/W�WO�!��t|{7�r����`z&��BQ{�'N��V-����Bwx{^�z�[��|��i)�c�r����'�,n�/�t�NL
�x|E����v���6���뙹�}o/\��@�m�Ǜs�|`	�y_�����V�G(m�A����r�z�M��ߓ��n��^�h��p���Љ#hr�?-�Z}���vS��9Ǝ �L�w`b�=��Q�Ϳ�O�B"-f��Y]t��#��|�1&�
�W��bv������D�l�; '�Y��N��r�WD��"jɖCڽoG�������dZM�7��-�/�*u�IͿl����J�4�|}|劭�qB��,5=<�X;m����,Z@ ��E'�5@�㏗��Z�T�>�_�Eoo����)tnGc#������6�G�,��d	L�e�⤍;�ɩ�r+�pu���8��.;��Q�6��������oq,� Y��,g��[�Ҕk��6;�\n-3�G'�.��������.��'�8�2�%Z���*-�5��$� $��?�l��ij���n�^�ۿ,=7C�x|�8��(�dJ�`��P@kx�%Y��<9�]_fC�TC�=���,o��n��Ə~f��D���to|���z)G��Bȣd1+9�ZR�w�,����k��{㷛1æ䕤����1?�,�n4u�淶;��a�/���00���I뤐Ũ�}g����OK��pC�:"��9���YwXu�J���gڭ���@pI1�d˂Q"�]N'(GܻF��G�1�����ܤ���n���E�H8a),_�L	�h�v�v7�7��e���=�(拾���
�
^� F�������	�3@ʟ�Vs���+�I�o�ƸJȨ��g4�d��q?<��#��P���,YdL�}ns���`'�x.���ی�q��x?܎�q�tʹ0C"C؄x�GgUd*&��r��/�{����1��/�?	/7���a=2R��\bkw4F�%Ћ�%.t��d�ǿ�m�����sW�F�/�/�����3�j�d��J6��M���{��#�b�O
��)m6]��U����ה�_�T�w�]��$���6h�,U��>袗��(��ø�v�o��#��m���{�}[{����|7��l�l���oJ�lz���e��)n��@�����0������N�����lHr�Vi�A�b���AhK���1c� ������.�='�uNR�K��E��Խ\,�=������-�����n�&�)���� e�8)�Q�Y�/�I�&�����YE��)�d݂$�qr������p܊qL����[`|�-;{s�P}ϱ��j��f?d�8�~�r>5������F�_b���t���xy��) �Ѱ�I۶(N�s�0���s��y�e�ev{�"{,#>!WiI�Ɠ���\S���0�"��È��0��[|�^�6G����ZZ/S]MBC�B�x(�=Y�η��`Y�:��ԣ�d�:�5k�Ӿ�
I�{*{��9�W�s�ѲT� y.�H$�����9v���h
ik�����z`� ���ݰ��zVHAQS�G�ά[*;2׹�Sb}@��Y �JA�&K�� KϮ���.��q��dT�-e"��^fy��(v���x�
�.�^,kУ=_`��ǃ���ZK��|��^�"����͖`b'��:�-t��#��P"n[�|��n��Ao��6_�Y)|�-��x&��e*XYqJ�%:6�m?�q�ntN���O���޻!�В<n��<�j0�!f"�sB�̏�ؚK�S'��E����'}Ό]]~._?Qe�K����p.���}��v	�Ϝ�jn٫�L�dx��$Fk\�]֣z��O�:��du	��q`�+���f��i.r��#F�P�s���W]���@��� ��(���K`E~�2e��=����zw�~ؓ�rϮ�4e��w�{�G�4R���}@��*}� D���2�U
�(��������_a�������F��#/合�u��������w���vZCT+}���+:�)�(FT�v���Vj��׼��z76���.�0/�p�e�	^v�~�}�(dG4��W��n�W�kAܾ�K�^�����]D�����%Fm�Ow2c�i�Ɇ����.˟8jt���|a�]��-3�T{G89�F��{�q�mL6a`q�Y���C��P1�����������B���9ћػ�r����~�C�Xr�]ak>P�S/�cw3�&�A,���׃D���C��К)���4Wn����(F�L�K���w�d�����o�Ot�x��:�9(xM*���b�|�F|
n�ݯ(#��<]ɐ]�~�'�ۧe�ly���؟^��zVƾ~�]�]�+GO�Z��4X����5ԭMɳ�?�U4�X4�T'E��ū���[���D¢� B��#f��
MR�Ђχ�g�k�3j��$���u��3�*���X,�����:�n�<�^�/���_sřs���l��1��+y.0N���~sϻ?{��6�s�'�*3t�_P}=�{��\�4�6������Y�1�E>��|o��WcY^��kw�H�^�<�ܱ0�I_�bv��*��Vh֧2[w���q�|z���~d�}�c� ���2�|�Ǎ��а�Z{2���n*yN�#�*��p�1���k�A/6F�	CbmP��	�e�U��E��-�L5W~W6���ŧ��tXk$0~�<�ɻ�@�E%�pM3�yޥ�O�,r9,����RH��bNT�`��>�
�N`��"�8d�ɪŒRV�8������}����;~W06�o�9f�~��`̙��,?���Y��_�O�n� �Vr!9�>ik���������h��o����M���AA�W��ߊ�|�|�(Lb����e�<�~��y��3����꤈'��p�v�@�y��Q|=|I}΀^���f��Yzr��M�W@���[����pW\�Mw��_�u���=k�\��>��z�M��8���I��/�V��\�dʕV;L�WD��뀯��-N����'/�����P��2��.Vgg�{����������y\�?Z0(0�-]�J��k��?R�%��J+���t�@�J*�
��I�����>VI�&��z�ܶ�Ni8y�A[�EZ��[�͆��I�����#a�v<?ѱ(:OQ���>R�Xֺ
:�|"PpX�D�|+x
�6�u����߭��u�1'��g)O����&��L�aի�/>�x�	������=j�{���[��.mM�kN[���5��bT�֑�>]9j���	��72�+�^OK�Gw��iU����״;~���|��rV�X��6PHκx��oi+f[����;���c4%X�%�TZ[��z�h{-1����(I����]��z��<������*���cޏ����{��E����3�4��LE�?�k�0�P�PT��ȼ�8�y����:���L�ԉ�}eNѺX����m�X7O��(p���<!t��� 捶}��7a��;I�5!L������O��/�w�\KǕy ]�$hq8�ܠ�	s�s���.�xw�,T�D]���q�5��q��Z�j���8�kj��>���"�O��{�W���a��]�����Si�_�9��`.�w���4��a�i�����'�C�p����#yW�I� jJt�'{1�zH�}�;���ۦ�W���
��b�u0�j��Z9VQ.��";L�� E��9��� �F��b�$�S���#��v����\���^�A{��.DE̥���9�k8���r,���/S�>җ�"7�ŀV/���OƩ�G�]}ҏI�&�V������Q��x�y����������M��=�&�&%
%=D��jĩN��Fez�����C���^��� ����a�i{k�O��/���ҳ�����Hkj(�l��t�BR=^Z\��x{A�<�<f�X����E�~�������i�j�5��G�u�m���t�����Aפ�lL�Q$]��Cn��L�Ē�˓��f�hh*Fᴊ	��Z/~��T0>��>�`���43� �[f���9�����o���d��ɴH6��4�
���_��;/��G�_))�g�#�8�^i�܁��{v/�v��p3��\�j��gU"A_�h���x� �WT�Ôb�:f��{V��*��5�pO@��̌FF��K(Z��|��B�~50���Ϗ/�WXeInZr��\o��:��-b��5=&ٽ��U,��NK$�A��t�����=�����>"+��������$��۞?O�C��f�:߲h0� ���*+���aM]���)JL7�M�/,�^�B�����ah�<��dXř�&$-;Wt/�D�Zf=���VL����ATE�?��5�� ��F%���u�Ƞf-0eB�C'���qĠ��1o�U���>m�Uu�m���T^�c>�V���[��;_�B/#(B�#��e ���S����t�&2&.K^!
�	�4F���t��S�,tIZ�����/�>ǿ�ux��x*�:��͑�eVB����Y?p>���`QICL��ȿ�d���0?JB����v^��L���_ ζS��z&V��3=AA�����K6ne^�c
�yħ��`��&�i�������?~�w��۞�����@����Y([�:$�'q5#.,$�([#���WhI���4����Z�S�1���-�~��Q�~iնTvF�Ɇ���X�Z�?�mTi�'�9�zUB*��Q���$0H��}�O��b�>�Ճol�t�[���&�;k	�+wC��0���~�ȍ��]���n"�=8���9�k��~zu�
�/rHBB�f/�yŏx{&_?�Cz9|5<ξ����-]ұ������~�6�ua��_�����<��~9[p�3/�,�Q&r�nT�f/��O�J�vtcq�WX�PIjOsa7��B$:Q���	�fb�|RM�Nep°�h "�|^!���φ�5�΁ӏWHëŔPRb�5�$*F���]�XX�gY.刺�tό���߁�/�1��4�\���0�J�az���.-�t��@�T���;/�+�g��!nBI��w�&;}��G+�R��6�V�AkW���=�ybT���Zh�m�c�=�:>7hϧ���қ��w-�����������f�y����N���NK}�(_������[�e��:��d�#�Ù%����I��s�V�Ѡ90��$8e;L���ŤT������ų4�2׋R���6@ɿ�K�`�V��0uy3D�<����[>�?�˿��� Ҧp���1���/Bg[�P�c��8|�#�(W�(Wlk�gn��������a��jkE!��"��kV�U+���Z]N[���N�ڳ��L�����5k�[�����w14���AP�t�F#ن�s{Pȥ䤀4�b�A�����&+UԘ��/���1�?��~�0lS��[[Z�l��,�4�g)(ۅ�b]	� S�c�4���pF��^~����gEV�Ud3ZyhAm�
Y�����ˤ�vhtD
�9���1LLW09]C[Wn��xm�x���EKE�y���ǂ�=h�g�l�t����Z����`׮ݒF:12���iI�]�g�Εp�]w�9m�<���ڼ�֮FK!���c�l$���?�W�xS���왏�o�"^x�|���؀|6��ݝh��hV��ҁ�����;�/(�\�0��W\����W�x�i���O.y���Y7֩����o�kx�/����E�,�e����@�j�[z �F6�`�GVi[�c�\�I*�ƛo����|Pd��)���2Z( ���#�##<R�n��)���
�l�����=�]sq������������[���at�����8s�z�SZ8>��t����_�d�	~Y������>%��yҍvY~4��v�2,[�X K�6Ցh����cb|�<Q�_�V�+�o<�W�ǃ?���1�v�_Yi��|�v�b��E�t��W�1��jU�ӱ{��}�ۦ�c..�~5^{�-�|�MY#�;�z�a��X8�]-y)hf��}�{�����!	FF���M7ŶN|�����G�c�SeQtWG+�[[��3�]�"�},W�ވ�]'������s������3O�x߀���v9%�,Oa��n�,h����˾_�%����Y�rE䊝X�i^z{>G�,8�'�\C���?�`|��MK����|�������=zb͎g��֋/�|a�N�s�����8�TAm�$�YA�O�/M��ڄ�D�j)�T$�wB �����Ojq�teuZ�_ſ	�Z��ew�����iH�ZZ�P3'G��e,^C�^
#K��Xo�@l��F����6a��%x����F:�:����hPA��m�,\4��ޅG�!���.<��څ��!��2��9 �i9_�O���\���
hbm���0V._�L:���9�x Mw�������o�Ï=�g_z��E����2k��V����w�����d����
����^��־�q���5߂[�?RT���F�qiOvf�\Ŭ�r��Q��ts��4\:�h��@�&�����{���U��߀4aulX�_��V����]��G�P���c��6��=,�ۍ�6��� �/ǎ�at�����C���Ԭ�]���%��{��zZ,d�q��6�t��5��܎6d��VCG[��
:z��E�zfؘ�p1���z|�/�����nK��`��f�CwG	^�.u/4l,>価����{||U��7ތ��'�Qa1#�kס-o��1=�z����% ��!�C���Jڂ�T6mފ���Y|�[���}!���8��7�m�<�[s�U&0���̕@��YKr|`=���)O&߂�>^~e'^�ut�w`ޜLN�!K�4��9r�����&�d.O�>:$�`x|}�CR���k��p�JO�N?��==8c�
��jǜ��D�^��Ꞙ���Q��rڽ�C:6�J�uhyl�����N��{�0�s�tI�S���իH����*�2�\o߾��烧'����[�؊�g���<��kh�t���`�#ij�:�Ҹ6�[��|�������C�g=LoW��;�l�=i���M��v9�@�l�/�RI��ƛn�"ۧ�{V���6��R)e��M����d]�+ӓ���P�����$�/�>q����{12:�ի�����CwO�-��M��U���1>1��Q���K?�|���7`dl�Uv���i�i�:,�;��))��hm�U&Q9vU�8"�@y�n��%X�z=zt�Ƨ1w�|����ڂ�Rmʺ*E��7��#�y�H�q�H?����yKq�����/��w����RBuziS��u����{t�r�(`��6�#��	%�{���]
;�Ž�?,,˪��T�z�I=���s��sϏ�\�#�acbjZ�ƺ�d�2<��/Pk����tt`bdՉ1�Y�i�?S��'�e��t����)a�'����F[�\,X��:�7���k����e�R�C̓��H����m[��?�|������5OP9>4�����?y��g��p�GR�_���<9�.��#\,�m�J~�H׽�{�L�/9�ɣ[<R̼[��!�|�(s�s�R�H�*j�Ϳ��d�8�G����\�9Tu�)i\9S^�����@̖��ף�����9}���m���Uk��H�
X���&�}x,��� ����+����3�|�=��wn>s�5���'���NKm6�R���A��/|7-���E-X0-E�����c�<�'N �714ڏK����t3����b�cp����T)�}��s�_}����a}�vZ������������?���D#L�dU�߽*��jX�7׊
��裡�h쇢���B�P����G��T5�ѫ�礫��U�*�5����CG
j7�^�[o���o~["Q����Жϡ=o��X�l�Ъ\K�~�w��c�6���RS2<1��>+&+5�����#�ˡ�����z�YH��5�������q�#���G���Obޒ��������⛘����s�����*9�a���%K�g�kё݆�@�TB��E���c}8x�n��W�
���?�Jj~Ų���>޽���m�*{�Ɠ��}���c�M7�il��uϔt�w���	��f��֮\���ע��L�����c#���k�E]߉19ڇ��a9F�ͷ���ߏC������aj|��Gk!��֢�2��W5#�� b|z
�#l��T�lN�_�q�H���:ZJ8w�V\x�'Q��YeF�?\�bK+ϻ����x��7Q�B��������g��tvI&�>��E��F�ɳ�	U�@��<��Z �:!��l8�PË���uSVV#z�
�|�mVa!֬X�/�v���kx��%�9���V�@k1-��F�w.��,^|�9�wvIj��w�X�+5u��ĥ�^&i!��\�b�og-�W,\(G�{:;�b>�����ǡ��q��1ԙ^�514:�����s����}P���Ն�"�ys���_�%��j�
���'��t��`��Rb<�̴�'��$�9"��u7����Զ�Z�Tj�����AK�$�k����G�O����{��:�;kt��tԛ�%K�7l�q�cc��@ ��R&�)_��IH� BB��`��c��;6��dU�w�^o�~���?w��f��kEke����9��������.hnm�P �Ҳ*L�:o����(%:Ȗ�C���=)4d�qhij'������#��a�FIy5���F��u��R\��C}}��c(+*BN�Ns�^��--ڇ�-ñJ݅F}�~FC$-�U���,�_h�X���>�0�����!k������EÅ:k�� �8"[�����0}�L�U�c�o!3l0�f���� ���"��GWV����g�B�ȸ>Bt���z�T�k��s;���)�2ιx.���m��gM��?�z��ǿ>�B�|C�<����;［������ c�7C�T�Df��8.�9[�A��'�hH8�>g�W�ȯ#DK��G,�iTd�1��F?�G><�d&FC,'	dN��!��T�A�柤(eh�śa��p6�*���IÄi�P9v<>>t�M�r�\�x�����}�(5J���7ި����o����]�
6��Sg��fc����*��l�v��W#++o����1k�L�>�H6������r!���K�b�J��]|��Dc) ��6���_X}�c������&������a}���W^�v�`���o��S��N�R�!'&We$<ld�7�_����s�����7�k2ٙ��_�,	��3]XapF�/:�h-��&�P���[�ē�G
��
��y�9��c|u%��Z�:K��v���ձ ����kn\��]'_ްQ�7uY'*�I���4/�̛%��g���%�i��������Q9v�_{3~��_���C�h⸱)N��Dc�J1g�L \�k@]]�
*I�23D�oiA]S+n�㋸�օ�^y%e�"�Ѭ�mK��لٓ'���Vp��)�)��vu�����n�c�*Sg����W�O�YcL�˼����Κ�+V,EwG�<A�ۚ%Kg�t���؏#GO��B#<�������7�ęS��AN��Ic�aWW�b���Rc]�ج1ͮ4���ڌں�]��r���**��vQd�y3f���oD^���Z��F�����7S��{�~��o@4aǵkoƮ��p��)�;V���a��Es���FoW;���9{
;w�Fvn���N�=��/��%�C嘉�Gbص� �	�l�Ɠ09�(k�AC�"Iw�y>�`7v���:�I�jP]Y���t8,����U+�SO<���r)�N�;����74j�B����oU�B��h����B4��� "	s�I�;{�a-
H�Y{�^�qr����ڱp�e�=w!�o�h8�L8{�SI~sr���Cs��E2]�g�Un^���%?�{z%�����$q���19��-(-����nJ�`�j�J��lvYlQ��3؇ӵ'q��q44w /f�]���ǰ?�Ü�<wX�������bѼ9x�-24�3�����ֆ�A?�ۺPTR��V߈}aﾏQ^^�1[oW'r�Ӥ �Lw����~�n:t@�;�V^�c�?��ۅ���D���/�Ǜ���!*Tc�����DA^�P*;W-_���b����Y]ظ����wpH��ӧ���[�ynW��/��iJAUD���JQYV
o��P"�b��Szu�������3f�Йz|Rۄ�ͅ��{z���O.�3�M�.���o���K�ϥP9}������͛޺~��ݩ����h1���
��%ͩB,�*2(-���n�L���#���3DSe"���|8�O�V;�B�FL�8�T��%����ڙ��$ӈ�~�I�b�,`����xv_8��͎��SQ=n��.4������˖�xJ��-�����b'��ԙ3شi3�/���׭�FGRq_������5::t�l���a5rr3��;o�bK���LY�|%�8~��ߢ���-]�y�� +7�݃�h�Q||����)z�ۯ�������������/z���_k����֛	[�N�����9{��o����GL���*N���d���)��wD�X��>�s�,ژ�M2��=���2�3����!��d�D0m�X�q��x��g�P_/���e%�,�%���f��<-����h׆[w�Y��<�	N��+6a�-�����+���� pڒ��Ge�a�*|��_BkC;�w��!�@|�$��<_zq�\-j�M��V�׿�::�1y����8�qd���溫q٢�8�I�
��]=��8Ӽ��"*Tں����Ĺ��������xX��C��PZ��Q��w�����;sVخ]�P{��Whbgw?.vtc��%�v�Z<�ӟ�9u�D�d��0g�T|�֛��ބ���#~�كCú��~m�$�vv�jF~�-w`���ط�c9����;�}lU�s������0�׍����s�kSk8|���0��c��$���oP�Ã�78���\ܼz5n\}�<&(�n�='�,7�@�z�o۵'O�Ů���09q�_������ZL�8^���fe�tx��\�G��o�Ǹ���]b��[X(�PIe5A���#��HZh�h��jx�P	��R5����L|�wb׶�x{�f��(��q�(U ���tz�Q^T(�ɮ;��6��T׶�PJ��8�[{�Mhn�(�ryi�����ɿ�hT�L�
�QQQ&n	����.�9sF�*�1��|��]r�r̙7Ͽ�
�sr����,n�()%��WfL����<)(��{��q�����������̂E��.~��^n��MM��l����W]���7V,[���Ŗ6����|� N�9�����s���X�p)>�P�)G?�ߢ|;;�+�a��2,Y8Ə���>�̗_/��(���=8{���-�����虡�KSc*�KDX%A��	X~��ؿ�x8�_~9�;�����'q�EƼ5J%�V��YB��~�+����D`s�1����}L��̝=�hhn�؉��Qa�b����G�XW[2�\B_��JE�D9#�p)�H�hϙ�uzv������q3fa�����|Bv�� #��� "���_�-������]W��<���}��R�tw�
F�����о��Z")��V�XJ��L�fqm�LY�T�� t�W:pS%S��##����ađ���h�9#|�߉�9,%��$��&���Fß�oIN�{��Id�0�P�$7�f�T	Q�:c&L��#�p��"LV��Vh�����4� 9����c8u�f�U5U���+%��r��7����<��ؽ{?�?��f� :y�V��,�f̜�����ͯ���7ްK�LI��Ѿ#ؽ�#� ,A�+y������.�����g�ֳ�E���7;��j���t{s���a�FJ0>#Fx�,�w�H����/H��E6�$w�?40< �$� ,v�M�65�K���z@��.=t4���۴�cqǭ7�٧����'eO�^i�(�.)B�ׅ�S&��,��A�:qB�纺z#h-+�-mhn�F�p�n�}CA<����0�� ����&4etY!֮��-M�����������(���:L�:C��O�I�nUU��&9^�fin<q|fN��§��I�yGw�
 ��+r`w�N�>�{|H��/�,x���Z�#�i���C�W~@���T�رC�qʫy��8�/v��@B�w��������Rܙ�cj�D�d�v��s@�&e�]t
M��{Pd�Չ57;>؃={�`��92z�"j���Q�uIy%� ��Nn�3;V:�rԒ�I�U�\-��4���&�`Yq�\�W,%�ӎh��A������;x��z�Q[�wz��:[�ۅ���^����`/�^:9�����jt��Ԥ�J�8�������Ā/���J�Cx�GEE�M0��)�$�[L0��"_S�t�}��Py��ER����1�(��G���"��1��s"���J�ذA|渉�j��V�Z���Vlݾe��ƛŁ[�h��љS'sz�!    IDAT��ڌ��̔��L�}?X���4m�,�_����o*hK
��v�E�7ӧN�3Ľ���[#&��������S�<�Sٹ��3o�ȝ�Ν���ۍ��v��*�5R2C+�H`��^Y=Zc�Ռ�u��с���܆�qXt�ex�N�1�y��IH}��&�cCvf��aL?Q�<,�(�o�؎ӵuU\�n^�m����={5�)+-F}]-�
�t�L�>���Bmm-�����Tx����b�lOd깿=���RT׌Ec��a��	Hs8t��e8I��H`��C���ޅ�m��0cƍ��7^��l��ѣ5�@S}���c�*�,+ށ��t�F���k(��i��g�f�L�9t��6 �� fu ����/�u�e�����wO�~�������=�+?��*==���H����V���z��F�|�p,L�rA��0'��=��#gф�,��z���&��Hj�%a(A�s�-{*	�b7�J�e@�2;p9��e�Y��P�yV�.Ư�)C�a,F�4�2�y@^N�-R0�o���0n�d��p��L��&J���Ts��℣���~�K���%���ة����Q��ÌI	Y()&>�����o��h.��n2":͠��а_�D,F,8�\���՗�}�w^��s�l;�W��K���b���~���ʃ��������b�v����@�T!i������9#6[M*�xm��h%H�5�HK��i�j"�kw E�>$#>�b~L?_�}����P{�V�v��Jd{�R�T�i>����P?�����%�+�On^>��(�z��7��_���><�`�:]W��$/K�����]ڈ�H	�K�j��y�p{������;~<V]}���Oj���:u�T���#�㶠���YY.O���ԁ��o�@��.���Wp��EP�^��ڮ'cA,�=}]�h!*1< �M�>>��4|�8MJ�=k�B\u����SPZ<JV�4��檕H��q��c8rx��S������/�@ZF���]�L���ؼ�l}�=u�<(�j�b��Y�h��űÇ�t#�-ˀ� �)tw��Ar%P0|eY��ˉO�c�	�=c�����^�>�\s٤�0����2)�!E��0�
�q��u���V>z�&MBQq!�ښ1g�d梧��uM"v���ˣ)7�0�d(_^����c0�b��)��%��6LR�6&�BΘ��Շ��wc��*J�J��Q��1�	�� :Z��u� ��6n2##3GM�0��x�a�����QӦM��9�ߋ�ӧ(����ŋ�:��Y:����#ׇ~R����Hye�.���_��+*����Q#+T�\li��L��j�RlfW1M��9��8u�F?�;��K���:�1���.��h�p��!�+N�WV���S��ޞL�23��ǆ�6���_�"�V"y�Y�c���Dks���\Os�����U���Ҋ����Ҙ띭;���}�n���א$U*�؀���5���"�cܸ���0r��x�D�!J����S������ō$r_QV�t��Σ��ɔ�,#$�5�T\�`(*^�B5cƢlt%^z�e=���4����я��ٓ��+&��v~�VDS?Fз'3��,TN���G�����H:3 ������\D�%Ȱ�ߝWS�՟=�Θ��}.�JC[�8����`4��7'N�P�'I�e�x�*��Hq@Ă����k��J�ŅD ɴ�!+��p��*�$��TT}*��P��%�9odkpOB�ܰ�m���5%���z��U�LRUp��b��s.F���xw�.�75#�rr��6g�t��ƕ��o,h�*l6��>�/%����;!::$�C30�8u�5�D6��n$&b�	�����N�[�P��$#�� ?����S���{��se���Ced�>���ط����^��q���Δ\~dn�#cr����m�g7ւr�}��h��c����i�ٸ��`hg�E��R�ܕdR�F	5��H���0��AL���]w܉?���2��}*-.��"/+K�خ�f�sScac��6l�nm޾` ݽ�����G����><�ח`w�ɿ���;�C�0#���2�s0����l��3B��뷳�Y�y���[��O~���N��Uנft��	�eE��8~T�5�[�d��J�!Ԇ��>�/hnm�O�3!�ӦO9����+Fi��o��ɝ�}6X@��OJ�@�y��Ÿ��k��_�F�Q�˗-EKk3��Tb��Y8{�S=�1b���;t/Y`���ӆ�
�G�Z��kx���������ϙ5m�-�0c�dt47��ȘmX��z�Đ��o��,]�L2ܝ;w`��i���O�Bks}�a;r�ϝAOW7"��CtEVVP�O�=�C�f�T�y׽x��p��	e"�����H��*����PT�[";ܫ����t 37�x��'iķc���i2�A��iu�F�%��8������C=������?ցH�v���):<v+��aXV��?4,�k�l�����&&�:��㮻U����?�u�7���ٓ'1��)��Iq422����[ ΍����"��U��ï�{�a��0Y�Y�p�-��[��x\R4
A?S�����qc�B3�2ssQXR�su����;w�x->ޏ�����PQR�����VL�*�q��q��app@*�h4��10n�$��~�ۺPVY��S��4��e��Ba����Ir�����F�6�N>7�����R����C�c�T��I��uJ\��Iϫ�q�P�ĳ����i�&cʤIN�V�������<y�^�B�y�)yV��t#��P0h�s,���)Eh(� g���-���Mo��=s�H�cjF#2�ǖ�7���%�E��e�V�ƢD��^��2�"9��A���8r�,����0��Bx��F�H��U�L_�ȯ����p�b���/m�ꪱX3~�HZ���Є������Ȃ��=�V�V�3�}<x��K�*{\U��,��L{iLuˈ���>R0$Ȧ� 'G�8o%�RQ��֎��~�Y�o<�hE�#�՘V��E�
ƚg核�D�jw!#'_�f�ϯ_��u$/�b"�
OdWa8�2��ຐ�B��v�J��� ���4D7�bBE�D\��P��ɱ�ao���<����ͩXq"+�bI��bM���ǔ����paU��"O��'__~�\˿�_���d����[(���F�UT2n<�Q18KDQR�$Z[���@����3"���R�I�ӓ�Q«dFJ����>Q��`_#8ԋ	5�*T~���04P��V]]%RnOG��!4xJga��)����
�K �X��v|���K�ƿ��*�r��Zc����E}���̽	ɣ�K��E ��O�d�3N����=�܏�󿠣�S�r���1�u��!�����9;���%�Z��k��]:�~�QIM���?��ر_�x���>ڳM��!y�V�:MD#�AW��.qe8�X|��~͍x�OO������fbԨ̞9��Ϊ�'��h
)G�y-��������h��q�W�����iӛ�����-S����@Ow���$R����(d��2P��L�

���e:(�z�-̞9'M@p8�-o�����,�3���G,���������q�͎1�&�kW��g�*�}(,X����O���M�v�Y�:0�=f����Gﭤ�TE6��&͜)2��{1�f�	�{�&u��+�y��ikp��_��x���=pQ��ǃi�:�
�I�^jF0RA��խ� wz�d��?� z���sω�C.C%9R���[:p�q�B��M$�������WA��_�Q���5��/�_��_��Ӌ�3�b�i�m}o�R��z:P^R���L�Fd���O}��_555�Z��
��8���ګ�S�q�zX��=��x���ȼ�m�c�N��OɁa ���q"���"t��"�9xH�F� Y���?��+
up��H	0��7���_{�w���qɢ��Q`_:j��)Q%ؠwQ��R���X�JN�����U,�i]�l������L�\��.�
�M:��xҌ������K�s;w�R8��Y�g�l��*ć*�ې(��S�a��i�Y�U���� �=n2N�5�ȉ�HX��{&�R�g�����n��?��䑟}����ȕ�Ӻ�s)T꺺�CA�/2rr�c)4��&U��F���a��f���%�hn��U]݈����
�V��2dl��6g�E����E=ҽ���n�����3'�Q
�G���I�d �a�qKP����[�'2�2w��������]�9�4Qڦ{���a�������RV�	&�r�bŝBR���"�����8̓8����#�G.d��8�$��P0^3�3M��UC�p�B(�q�rٜo|��e�O���[N5��-������2Y�Ī�^�=�ڀ��!��'oE�L�,�[�X�2���B����/�H�L$7�*��l(���1�(fب!U���2#�K�?�x0 D2~z��{���<��-)��(Ǝ�уOG���R"�Im���G
���6���1�����g�
�ͩ�"�bȇή��%9#���H�Thу�8��%�,�w܁��q�;}�}�}())CM�X�Dy�$�4f3˙��ݍ����b�ז���o~C����Fff&��"^DC�i�}�"��L��ݡ"�C��S��zN�2��q7~�ӟ�V���@sf��z;~��\\ٙ�~��xx3q���g��������?�	���6��Eꢼ�,^���8x�c9�RL��쬌��v���M[<fx)Q-t������O~�{�`�<TW�`���8v��b>+��4�$Z��_��Tl�N������[���W��ヒ�WTTaѢhim��C�[izf.��򅆴�4)[���>�,�vf�[ �ۮ=�%�%���$�P"�I�O"�x��K�|�n����=f��Sk��p�t�mmQ���1�f�~�ṽ�I�JB6�p������ڦ��"H��DYi�H����8u��"���X�B�8%*̸6l|��5������~�����0y�r�>q�/F�!C$��L�,��!�I��`��I�~��I����-*�ȵ��H\(0�͌�4'*�������5G�7zˤ{�]Y.���q�=����p�gfd�:456�~�>���>�{�G���OE����!�=���V������gh�`��p�0�d����X��u`Tl���~�z�jq`��܋F��)^�=�b٬	�|���ddzT��	��EE���g� ���B�"���T@<ӊ�J���$��EfF��x|~�.���L���8��&r��+Ë�ʱ8Wׂ��M��ڀ�~�4Ձ&?��[g��ȯZ����ǿ.�ʑ��ꓵ	������E�t�����1iC׌��76�&$���9��a�6�i1�踸U��z=nB\��b�����a.?��AΟ�ύ,�������x)��Aɶ$e��#+��2����Zm�
�N����b���kh�n��cDF>�>9ʣ�A-�Vz���ʐa��eQFֶ�qX%�e�O)�q��aac���#3�E'�>$�C�F�M����_�i�����6/�d2i��׶/~��ÏE-�yC!��o0l"Bs#���=�UcqJ�5B�O��!YWh�]HZ>�����@mp�Bk�W`��`8���dMο�[����t���^��H`�fN�=_���q��I8�.��@���G� �{z��������]������������?=#ؽoxP����C�ʃa<�fv�<��ja�c�k��Ӆ+V���nƏ~���ɫ��,���� !1[�F��^�W��I�$�B����(��O�P���xf��[4�@Nn��98�CVV|��T��I�j�4!��A9#+�ĵ�߀���w�����j���<!�4Vd��"Ðό(?320dO�QZT��{/��
���]|�xѣ+�Q�����xeD6�,�L��`7����Ӝ^�]X����/	9��%�e
m��q��1�K_&����TɎ��������~�LqL�4�<�5<���8v�Sجn�2�?�s2Q__+;��|�G��#��ܰ�ܳu��Zs�M2wۺs��>C��x��K��Zq�;��N��i#N�8�ul1Ӊ֬k�MLr�����'CA�3�X��Z���wߥQ���_���Q�Ak���� ���1d�.}���t+�1C�2fWq�Y8>��^���?U(e��̬2Cd�X$�B��H_d�y�Li��\(�����ӽ��w�/�Z^x�ex�3�}��
{��a���ix`N�"���͔s�̹�0i��%444#3+G�5��J<W�:�	��Mz=_PH��4�X͑`��
�Y�7�.U�)��(aȫ�znV���`~Ѹ��WD?�C�]��s�L	_x���@DS>�6�I{t4�G�J�P��?�w*{�	��糵|�r�f���^��.�!&�ɦq���3�W�1�����As:��pyţPY3�-�8Wۀp,�B��4.u9����O��M�,|�w_����(D����\
���c��}藡�}�@(n��7�&Vnұ�
�m"���2e�΅�F�-U<�Y�pG�<���0L�F����u��(s�Hu5k���-�Q�H�K2FWI�36UqR)�"�Ң<iH]�1��� C�
b(v3G9�B\J��	c��
�(�ń!j����Vua#��~��p!Cf�×.Fj������	Fsmr}XUH�vj��k���0#�eB��J3Gw߰�~}���6T�}'ƽ����k�ά��Ń@��E���swI"� 4��N�`w�1��bU��*N�� �P��,`y�5���@4ʰ0�>"1L 5\m���Ӥ��4�$���b�R�̙���2~���h�����Ơ�].c��uX����.�t�e�=/���5�����&U��W^�Ң�YY���Ƨ�U(��hm�,�̀�l�G
�P���ߎk��
�?�8N�<i�	�����hS%r��C~�23�޸.<�ƦN��}�{R%��oUw��"R�8L�%b
t���5�T�� L�|	�n�׬^+r�O�k�<}&�1��;D��@�a�h0xox�qq�ޯ��>����;[�ap�/��p16ց�HlV�l�>1�HhV[B�1���rr1��<���"��ϙ����E�ǌ�HX�
�	�}�<i��	�	�ˎ9f	�����{��q���de!++�'ǆ�/c�N��P%&%O��I��k֊��s�GH�,�#8j`����ϯ�hc0 D�ګ��X��}����q�>�Tlq�0"�ׇ��L~� ��ĭ����/��_������u?����i��!��H�+9vШ�E��c��X�j�B:(����+������6�L>�d�Q������"�3����p�����x�ٿ�(爜h=A��촛	�W��J~L�~�.�=��f��q�Uנ�j6ozJ���=�>/��J&'^o�}V��d6��4�!x.��w�ҥX��<xP�I��iX���4YG�G�Bz���1|�Y(F1~�X�|�:!�[�~M��ą�Z�]ex���"���(����1�9�R�%M�נ�|��Ų�س�C)Ҹ�4rJ�ޓG4�F,�g%I��)�7J�5���ӑSR,O��n�a!
h�K��N��g����;�O�(��?T�r�k������,fI[569�B���� ��b#/�2F1�t��<���Xᏸ�*��
Ƙ�9vhX.첢��@�oaE��5�h�E��e���7#��LG�4�R�J��z�u0;�Ge�|ΨVY����,���s-IR.1q���ϲ`�K��HMm�|��Y��gu��tb|ﲊ���	CZM�J�;srbX�=�������9EV��P?z:�:Ks6���~{�������7������ֵ�/�|) ׸����&�RI�����8]�ㆽ}*��0d���l��}02}L��N�9YF���8R�E��dO�Q�{�ڌ    IDATp7n|йɦ�y�Nx]�6�	�U�������R�~�zyh��P}��y��QaD4���$os���|�Q8d�7��o��]^&|��� 7"�|Z9���RN�t=6�T�������/b���2�{ꩧ4��}4Tq�&�XA�3�!4��3
��ȫ�^�K.�T���o`ӦMB���w9l�e����e�|���j�O;o�`�6�K.]��J+?>pT��
E#'��h,,�X,�wr�2Q�랖��ѥ���-F]}�~�}>|T���ݢ�`�r�F���H��Qd��{1m�t���]���N����p 3Ã��n�1�o�y��T���3�e\�Ϟ��S'�b{����Ga^�:����
s��k%$I��Z��e���4:a�T�}t�T�"N7"ɤ�gcݙ���s�p���:�N}����T�����d^_�ǹ��L���bQA,�b�?��,�7;��$	���{2��z3�F��努F�H���g�� ˜�5s�hU��p�%zި:~�S��wÛ��H8��P����P�c��H���HZ$B�5U\�P�0G�Ѩ��O����E�
�|<��OYR���2-��TP&�Z0E���4����ƅ�Qs�E�oY��ˇ#�h��<Idgd�`
�B�9Ng�Ȝ���j̙3G�hX�ݼ&�]�Z��EeFB��iCQQ!��2?����,��Ԏ)S&���sˌ�� ,@ӿg�4�'H'm$y���:��نH�o�NNf�8���G�'&�,�<��>Ξ;��F�e�_�n�:�(=�7<'�UQ��q�##��,4�w��B��!ܷ�3X���
�9!DeBE�?�r�+T��[�6y���g׫��_�j�`3P���$�bY�UI����b�����U��њ��4��|�9�#A4��h-vƄ݀i9z1�Cl#`�"�Ag�Î����V�VXL6�,F��Q��0��#'�]�kV��i@��F��:�mIL�c�)�7�/%l�?uf|������*/)���x�(�!�w�Ν6��u�^���5��be�G��z˵O��H�&��r���`nOB��,z`�2Y2�׎���v�i�d�(�X��!d�k�O� G}z�z����5�h�
m�̝!d��� ;+����h2��$-$焛!��W�Z��^�p�zc��C�i�!����.^*�HT�
�D�/?Q�$�ϝ)�S^k���D�3"��MU����3����z3�e�������r!%�ѫ���IA�2�_�2HvQ�<�/��s6͑
�;n�e�p:�8u�
��/_������B��~��!� ?����+rywW��{�.'���T��DN���NL�:[�q{w�!��-r0u�m���Lo��|"���t,ٹY�f��	t��Ø2m�L����~�h�2��]2莳x>#�U0=�b��Q�I���;�L6n~=����;�^M$�Ds7tK��ܖL"'�����Aw� 
����Pu�M�����N�Ï��D����A�f(3��"o��`N�ɂ�,�>C!��h]@b4y�b�9���HZ�2=s��h�S�d�vl�H�es��r]:P�	c���#C/���z0��(7S��$ɦy��	#o�C^c>7�o�.��o�Y��Lu�XQYQ������+��5
S"��[H.-���g�����ʊ��kVv>��3H�_\H���DU�/F����+b����,?��[�nAFN6�p���Q�΂-+݅��^}}���1>U+�@i���!�ݙn�OK0Ň{�)fd�ʕ�1u��lr����f�Yb��t��y��Gৌ;n�����8r�(�޲����(�|)�i:3#�-m��ͧ�~�F�l�X ��`Q�Q>I�n|M�m劫�iry�*�X�RD�q��$])�ED������	��|4�#��k��3N�d#�5)NO��C��)�7z0��
�Q�ؤ7� N�7����@�$��c�B�I��/���6uL�?G�pgh�w�$�H�*�+@��U�<&%3�4(D��WJ�,����N"��X<�{'�2������##vΚ�X�kd~�x�r$g�IX$��ae�P),�;�LBl�I�8�g�iL�}̞��3QʚS# �"�ܬ�	m�92�����O���pUF����:���"c�m��&,I��wn��Ł�4/6��18 �>�.�:�;j�s��Z�l��-��Ud
����O�ynǧ�_{���7�\7;ǆM6ON�6�Y�=���Ε,t��q1!;Ia��3gڼ�D��s���<B�`G�8�^'�Bv��sc��8��[$�N*�>Y�����܀�Eb���u�8y�O���,���{�L��Ka��}��Hz�81�P�Z�TLP�y�WJ6y��1�ڙ~�0$�,Rɓ�{��B��i����ұ}�6�����Z�4��ر㵶���M�H@Nv�|QJ�a'Y�h �=���S8u����!ݛ��1�1w�,�C���n��y���B�Ν����/v�'���<���!z�߇'�z��_X�ʪjd(������E��E�T���p�z�E~䌟Nʴ�?v�89��ͨmhA2a�رQV\.��\�gO��9��q�"�����r
D����7Ѓ�nqK���_���]⊑(8v�
�xL�ű�0�WWaْER|!3��'���;[w���BS+���՟��Ȩ"�j� ͙���r���w����ݼV�$��D�g>r�o~S�,T߰KolkC[W�d�,T�"p�I� ���H�)ԌHg�Y3؏k��/m1l��G�ˋ�'FG����Ub����i���G�3�?����*��Cq�l�Gr݊�r\q���/��/�"W^�ǣ�&M�ZZ��vy��p�M� ���i�ի�`Ų�(�qQ0���#2j�7����¹�H��fd+Գ��� ��Rx+���(��?ЃXhX�%�f͒l��=��I��H�U2iS��~�Tr����df�)a��c��r\}�rL�:NYMv;p�L^}N�<#/#�H�h���JuI�=t�6�MA�zx�T�I�b�T���L���6~I�6ا���1�[\'<HqHR�<�E���Xs͕���ȇ���#�r�x3r�?�OM)&b��� _gR�DHG2�fM���3g��W(S���g�~�ojR����'���[{�9J��g#�gG���>m\�ÿ�GR�j�ڸ��O�b��C�i·S�
�g��O�aM!(�#4��\�d�ܖ���!��r�S��<)8g�@n����`a�Y�1�1XF��D���NFc���D�b�:$ϟ!wE
��r�!J��V�q��18�$��A�0":�W�`�s�����*ȓB��2�e���1U�C#�g��b�Jx*�2��k��ͱ*�T:�����@pxHs��d,��Z��=��N�~e��'��)�W�c<i�/_��������{0^�'*���I��tD��R�BX3)$��e2�@4�\�a�HD��� И�f1� ���-h�p�g$'�3ov���y���!?3�e�
���h��2;nBἁ,@yŹ�?� :^���1��֩�N�F�:��h���%Rl2�%�,��iSE$����/<�����Q�UH o)ݼ�~���/�.��W��\��m�V��ʕ+Q^V���<|'>��c�L­7߂�</B�a�ٙy�A�3Ͼ�c�k�rg#M�1�!��EF��.[��nY�u�ʆ�@i^�=n]w3j��18�/U?3�b6��	��|"C1fS#[RYIW�\���^���eϟ���a������`w����M��E����<�hREZ$��YSq�7��|��mx�ߟ��D{���!C0���߭B��]{���m;�g�ʠ��! �LBC}�j�2|��Q�����qT2�
��Ճ��~�w��` ���$�Ȑa��6�œÒH����W㞻��΋�hjlL^VV�D�?<�'I�y����_�t���0��f!��h�(bSck�k�?8=#��χۭ��+scH���
\�`.l1���i�a߁�x��*�R�CA�6e�n�I�KV��/X�� �.�.Ę1c���x��?��su�h�,�'�U�5�9d�iܖ�S<���||��b���0'���dWñg�q��7O���V#6�n�s� 2�34�e��%��Ú�5I�y�.+V�X�믿^Fz?�鯰u�.ؙ�D�>i7� �v��̮s�#_>��u��I��݈�n����uFT���j��u�؄��>\l�4|h��%q��b&���,,(�Ș�#�)��j�c�R5ʉ@L{�]�� u�^��1�!�9�Ԙf��	��u2�۾u�
(>��	I�2�*tIj���<,��_�ԑ?�杅ٵW��̉�p�yK~2s�QV^����w�D�?{^!zD���ӌ�{��)CJ�:5���1�������$O>�1P��{�<q\;��}1jR�"� ��C(<5�>6�)?�牶��i�a�tC�!_�hL�.K@
L����0��(��0?H����5�	Ê��>"!�ф���2{K��ʯ!E���*b�)�<��X	R�aG2b���A�x��+5��P��FR�ȗ�]��7�d��ѓ~�ȋ�Y��Ò�*dz��JD�._��� �C��[#`���r%1Ge�iO6f�YN���=��xiaZ�7-=����㉤�ˇ��n{}�?��B����؝�#fZ�n-��q�f�C�IjuI������P�B��߰��R8{�x�+Jt�&u���d�ӂ;�73C9?����]�JF�"�Q�<s�ܼ����g%/����q$�Cؔ��p�ۿ����T9<0���"���dRI ��j
���zmP6�*�#1�U+�c��yxg�f4�4���d�"t�taǮ]R-�K�.o�g9�t�ri�R}"
�x����Nֿ�,�n�S�L�'�+/o�L�f��˰��p��C���mp{lX�d	�_�/��&6��T_�u��2~!��'nY�W��J|����"v��-C8Z�/Z0_����?�����W�¶���s/(���c�7]3r��T��_{�fM���g�˟�T�pD3�/��=p?2rr�_�/���/�`Ζ�M4�r�S���}w �ٓ��̟�A(A~^!��o����7����Eey�ΟOz6��59yV�����N!�H�o�a�x���`�v����۵����y��{������	���U�Q�!ۨ~�$��f��|W,��?=��[�GgG/.]�L�z�/x�n�,v)}`��������9��!�=Ո��7�,��d"!�G5R�(\6�=6�C�Nsb��YSY�9�bl���=���Ǐ~�+t�*���S���
}>[)������0JF���֪$I��#��hi�/�@�pC��^o����cXe��8���̩c��o=����'O(A�����6�<ӈ3u��R�Qڱ�f�/�Wɦ�Ȏ՜D�ǎ�P?�=V,[�7ݸ���~�ۧ�ʫ��Mf����B0�0|��&�њ�����H��N[_}�˘8�_}�Μ�A�7��mqZ~��ߪ 'i���*=C�wݚ�jD{���k����P.oT��>��N����`( ��G�T#��c
�gı��^�89�N\y�2,Y� =�]x��g�z�	�ح.9&{3s`���,j��HHX�3&���1Uz-�͂mﾃ��N9⮺�jXN����h��Àَ��	3<�Ē����?�j�-��
�%ҿs�Ģ���?�������7���߆���!x�݃~��!���Q��2�9�s��ч�r���k&t��n� �?���%���P�0��ե8()Uψr����S�#�*G%\d�D��,��8�~�P�"'�x*Y�1d���g�ܚ�&इY�LD��i�
 ���͂����THDI�5�9q,��%�Q�(�I�y�ӝ�]Y��d��V���x�H�p m���s�ŎE*"�\L� 7'��3ේ�}vs��w�4��V�=ǭ�7=�4'͎�xk�۽1J�\%�$�/�C�H#���!;;yy�rq��ƈ�`f'�aA�o��u������.�	a����AT�Q��(͎�o ���{n��*�|��lø15z�ׯ�E�r����uUUU��W�«��*�%B�*z�pὼ��$#���\�[��f���7K�
�D�[��2\�x���G������9�C~����G<��}��A�۷W�-�}����f�=�0�N�"�ß�xJ������Gk�S�NiC���EUE)z{/��Ҳ,��R9������ڦm'h�oo# '���2q<n�������Wq���ɳ����DsS�/6�q���a���i������!��*囜��%��zl�5c2��ve������6p���Q%���[q����?��N!���6����i�r�p�%�p��7����w��ba����DvN�G�����/߫b�g�GCk��a Y�#zq�l������֠�����H�s/�����k���WO��/�~I�M�v�,l ǅ��!�f�p�7b�u�0�׉�{�����.]���\������g�	3�:��MH�H�7�*���}`x��f�9H��ʆ�{�gw`�$	i ��m�#�iAɨB����QZ5;w�ǳ/�Gg� �N�2�F8}�(��3��cBi��|���T����Ml߹�mr(&���d|�í"��k�ʜ�����Ӥqex�_��A_g+�KKa�{�ӉS�q��8[ׂ�5��C���u/=Z(���@���S"�z__��6deР��1���^Ć��D4nB��0,�t����Z�"�r�7�Y��t���LQ?�Jr��"���(������14���ϸ�։@(&g��R�]�s�WsH�䳹����\1 l���9z�w�B��Nq�LV��s����c8YKȑ��O%���y���!L��·��54]h�sϳ!5I�K��8�M٠&��x,*�]���@�?V������[oA�?�-�7	�垷憛��_|u�_���ف@ҊD�{�](6ME�#go��Mq���9oZ��G��?��W��#�ꋻ���4?���>:�FD��Q��5mͣ�%/����SB�l�C�61Z��$����4%#U��Lq�F�^'숉e��I�WR�!)�%'��gD����CVRa�lX���<�#���!?������f=���ev*Y�eH�����{�|<���
�Fȳ�������{���z�.��Mά�Zș �����e�b�*���<�/#^���G�A>� 	 ̱�5���X(�GVK4a2'����js�L6���p;c��P8��6��2�b���c"	�i@w߈τQ\)�Q����IT����A�P��;����hH�)7�in<�н�Kw�������\�TD�-[���\���<���o�xQ��n[��{����Sb�/[�\�Y�}�pO?����J+��X����x��?��R����}�m��,�o~�3de�c��Ѻ���ցo|�0~�8>|L~&��(-)��/>��F�����BwO�6�4��-�����k�7�-��_y�ORXᡃ���ݡ���0k�^���*���E�/?�v��g���4��jI���"��\�ɿ�fL���Ç{�V���t��1�׮�5�^+��/�;�<uND��� t�"�0y����GQ~.��?+���5i��+��o��������NX�C��,Y���>�y��l�l<t�ݨ�;���H�L*�}�Q��V|�;ߔ����[��]d����x
�j/�#�p,.�[s9\8w��6,�3	� UA�]VD����{�'?�#�#Da�#�#yX�3�� ��o�˗�S�^�����l��L8w�x�i>v�8Ǵ6�I(��$�yA~��m6����0UqI�a�{����-�@    IDAT3̉��~�#A�9hz8s,��c�p���`���xo�<��F�v����b�ya�	�p��,"����rY�ŵ+q�ʥ��2k�N��j��ֻ�q�t-BI�"I�Lv�h���xf�$���.dg8�Ő���/�L�Pn8������ 37|x
O<�"�Ե��g��=4��dh�j�zGa7�㫖/�?=�2<��@��cGGw��)���ĩ����&�t{�Bc�"���l4�̢Hs��%���@A^|C�8~���o��!υꦯ=���ֿ�cG�@.ǘT���ۯ���Ŋ���k���X��u�jz�|"�Mc�IN�!��S�;,�	���:���}㑯���	�m݆ή!�q�]#)�� bq�q:�Mr]�er�;5",����������_��L��/�-�S�<���n[l&x/ɛ��Ԙ�W������ms�<�Ǉ���IO>x1P���}�����ۼ��II&9!o!�"�����MC�Լް"&
Ac�\:d�2�Aj0��}��!
)�%�"
�keD��
ƪ����Ⴉ�n�3��a2H�������۬t���d�F�a�iU*��0�3�U�}%[w~��a��,|����( �Ϣ�&�sBY��Q���1�:��I�B��r"��$0���(�Q�Є�	�b��_2Ww�*�O���zM2��b�è�"�G� DR(�fQH�,�$��y���B�)�#����#0"��3J+v������B�Ȅ�"C(�MG^f:����c5������IB�|��hݭ�cÆ����Z�.Y�u�܈�_��dݺu�;_�l��QE�1}��}���8K�-Gzf��֩�!A�7؅Gy �Y^��׿����p�u׈��;����߱z�M�Cx�gp��
��ηU�����L�(�s�>��F��;��%x���(�^NN�����`~�����a(qXN_�4ߙ3&���P�=��G?�=6��1���qI6&z�� 7ˍ�|7�/[��7n��-�ae.�A�6�5����5�����;í��n���T�ދ4E�� {C�h�DKL�є/��K��$&�X�R�^b�����( �H�vz���v3�;ׁ�?�W�#�y�`(��5ל�;�Q�lنG{�7lE6W��>��J]K��,4jk+q����ⷿ��|`��w�1{�������g5n۵�	���h��Bey%|�P�#�I�F㒋����kpۯ~E;H!K���2��_�*�3x~tݍ
���wᫍ[����,M�k��,�b&�D8�Ѓp�!�ѿWOĘl=l jj������u2�
�(;+d�ea�r��j	��г:��.?��<V��/�A4bԁ����y��˯!N ����9M� �~,xP��`�N�;坙5|�U�;��B.cE\W;B���R�L�0Ι��S���ח၇�cӖ��T[��d�5"|,��J�L���=���k.��'��E$e�O8�Ĳ����c39� r�&R7�I�+6�q�mJ%>�7.:��3kV.Ǉ�����+�F,^�_��'����"o�K9CL5&�Kd�q�O<�^4G�rpH�.��c�����#x�w��Ƒ�/��'%�6�g#�C�E���AE2 ��_�8֙R؍9Z�ο��w�d�r96���5���K�5��I�׻WOL�<�� b�I�䝼���8�sp��x�����o �UB*[D;��i��kߤ�%�ʤ�qϣT�h�6j�P����c�<�ؓhhj�	G?��`Һ�4�<?��8��*�9�ϗ�]�_�B�l�ۚ��/h�N���sg#QY����������R�螙�yf����"�\{�/��A���k/���?��o1|������W��Eg>:+S�VR���j�;<�xq9�ࡓjm��PI>+^ -�My�G,�ʑEC.��0��]r���S�pc���L״xݡ�+s6�!Id�)������v�]f�.�4;:�:{ĭ�5}$$	,�d�u��$[;��b��B�����x��H�r�u(?�G�%L"r�]rS�Ǫ\hq�	���w�uf�A��Ť.��*�N��kA#�Q��D5�%?2)�E����i�mu��*�+epF�Y��I��F�KD�
H�d��K�s�=.������lu��������,�!Z"b��H*!t�"DmUn��� �_��6)�p�q���ϱt�R\s�5صw�8+����l�w��;L�0��p5�-�
���5=j1��IRU=2w��N>�6O?�>_�%������qȤ	�ɭ7�����1!3�Ν��~�g{�tqD~{��ܩ�\z1��s�|��0s�t�����K(K&��r���Ua~���kA��[n�=�)Q�����.�5v$N;eV���>�P	�^t��W{�m�7�I�5��@�1��}�Y�#��W~3N:<0W�U<���)�'��c�
4��y�h�Rq��ʪ���S�2������t=��냟��*T�q���o��{�{a��c��ds���'���/���ô#'��]��?[�;{G�������ŝw�VεCǏ��յ}�_ކ� +����#�u��L�q�Q���iS�|�"|�l)z�T������g����m�/o��9�t�`�����Rfs�YU�´�"��n��O; _�؄��ˀl��0��qX�؛x��*��8|����9V`�o�
9sF��k7�1�y�N4�~%R�ٮ��+u�"F^W'N9�X\��0�5^y�<���ع�m���h�D���hy5e2�#��>g}z&q��W`�Ac寳b�*D�q���=p4n���hٗB�2�h�Cb09p��@6�`�dԇ>�9���"��|��={�~�0h��~�x��h��	%���:U �X!r
��LF1�_�r��àm��1���3�፷?�����;�D�%�m{*q
�o�b�Ql,��s��P�gG{s=�8|
���UB�8����e�]����{��ʕ_ꬢ���G9�#t:�J�ov"A��l�Q2\�W��.� o��O>�[:�U���!	��^�Z����0Z���gFY1+�ڳN���g��TG�<�M���R���B#;�3�t���^P�
+%~p�>�h�y*�_���Jq<dΙ=G$����۶���n�R\�1)y�LQ�� ¾|{~��^s�M߮��W)��P�϶��y��w~�+%�-Eʫ)%�|�_���I��}�5��q��U� ��X�fafi��7�\׌xʊ�W�D�C8FP�5tD�I>�\9�<�.�+�1H�cJ����<xHj���Y��(��X͒qI��Hq|U�7�Y���G��%�V���X1�;uW�ڸ��d���aX��wc+�؍Y�Ƣ�`e��m�<�Fb��#G�+%B�̢��3�=GVW���ha�c��֋yK?-�'VƌSWQrZBHh6EO3B#���,N��KgT�I��{m�8^-���%ˆHM�<��,TL��M���#�6��#�6�^}�}��{��}�\s�ՂD9S�=g�T3|��#����_����k��r܉'�`�8��Tf��[��^��
�A��`��Spם�LS(B�s��8e�	��]�c��ը��ƙg�-f���1}ƩHe
���$�����o_��;T��e߽T��駟��4�ꋟ�z�r;��ݝ�ևM��뮻
��Z�x���{����Ë.���:;�n��o����r�'��xh��xp�Sh#7)@� r鴒m��c�����`��jh�<�֭݀aÇ��߿#�R�ŗ�c��u�WK�~���#M��-%U���,��p�̓pک'��"��{O?������yɥ�b���X�v7��}o��!�D(T���������s�©����N,�7��>B������7c��	X��r�ٻK!r��-��৿�5�޾5���u��˝�"ƹg��4m�|��{��38t�T����_x�?�"�� :��� YV��� ����7�Dx�]t�9�p��H�֯��=j�hȹ�������iL�Q�OD����Q��5�g�e�S^V�=�U���2i�5�#o2�Ǩ�q�5Wa���x��O1o�l۾�bH�r8rb�_��7���7�y�sT��vN:~<>Y�K�.SAyƙ���r\�����eȱ�*1�3&2-ɘR�P-�cZr#��)kn��M����g���1�Q8����U���݁%�� U���D���q��߼��RQ� �Q����_�������,Y�҄��⣚��z�����R|DhYLq�7�OO����c���X��lߺ���´)a˖]����b��8o�̝;��>�D<���*9?U_�u{пW!��)�5������Ź�/���O�o�޼v��"Z^�X�;��VcIy:�p�$����1f�\}�w1tp�q��Owa�܅�U׀\ާ{�q��2��\3�D<y^�i��]�SO<GM�����^}+�銯����a뮽(2�!E0@�7�s�fs�s�@��|[ԗz��q�_��,߽��ﯸ��/�^c[�W}S� �$`ɐ��]wN���Ш�9�r�pFHdC>�0��dձ렣T5�tH�
ũ},�ǐ���E^���ȇ�iZ]{y1ޘ�Ȃ�ވ��`X�hP�\
&53��#$V��ɜ.R�a$;�`w%HRe��Y��}E�Y�[c��r��w���ӮFFBIĔѿ�*��r��#�qT�j$��xL��щ�0	�C��h
H$����ť'��"�	ݟB	�M��H�0{t3֣���aAj��̫σI������"�WJ�ힳS0��S���T`d�b�HXr�����X��j<��|��ZE2�u�9���99��x��g�n��p�	�,Y�Dv����SO?k֬�[Ｍ{G���[�"��'äI�1��#�ǻ� 5�f��L?Z�KMu�w�LD��Ͼ��O��K��}�w���hni�rŕ�a����헿��ܬY���Ԩ��z�J���'����+_�o�	C���>�v�7�y,X�(&:s��ƴ��d��Kk9b�����k�l�?��<��������U���W���{ n�=�,�x�Is�Ѹ��k��!�#���� �~n1�{p���|=��~�Gq�Ap��?���嚻3���܍w�}Wh��g����{�s���ߡ�>�B%�������Ӧ��W���૕{q�����-�p���p��נ��E�s
�nc��x����֙C)A*����-��N�������r����d����|�{�yu�mD�$O�szN���=��Mi����İ�}qݵWa��*p��.��5�/�S�>�=uM�'4�1���Zx��4ˎ����|���&0E�c�Qr�Nu��#*C2�V��y�����\���n��N���֤��Ze	u�l�JD�#j�a�^"г�"���)cq��.Ű!�����^��>�=��@0��/?�n�
^rJ�R�v��g5���pΙ���΁O�$C1#h�,��c�O`wC�Pl��d���{gqZ��|*��L�i[�P^���
'�|(���'��{�tps�H�?��K�i�鲎$����=Ѕç��\4#G֠*n������6fL?�n����S�Ǎ��~}1v�ɸ���a��0�x�L���6oۊk֠�!8{��x����� �#�2�P����H�A�(]x9��be��`Ɖ�k$�&T\<��K�ͰPd<��K�7�)Q5��X��4<`P��8�#0f�h$�!P���ux���ذ�k��Th$�?@�_�?�4O3C�s����E��F��f���E��R��~W�)�Rd��?�~����` �������H�b���BLF�?�K��9��#���k5�WJ�2_� 4�x���C_�����Or2�^Yy�L�6mވ��Rg �%L�e�������8R� ɽe�L9r��~�F⛽x��ױsoJ��S��1�W��ƓxJ�ZrY\�����c�&��q���"��SA	���K��C�	�[�TVZ)�pbWi�А"I|�C%�<C��J1�#��oh������kۃ�!&��@�uU�]�Gm�6
Xd$ ��-3���5�˛�stm�⨸�t�o�
�ׇ]�����j��w���{�\�����O������I���]n�_|1�{�i�[�Fp��SNà�ð��'D�>��3p��*����;ￇw�ÏT*�IO���S�`ޣh�<��
=zT#�����}0q�X�4W�u���xl�S"�6R�捛7)`-�M���?Y򙺪ٳg�_��Z��4�Z��,Y��d���`a٫O���}�}�!�4� 3�0T���\� �۵�6aѲO���E��u�5����C�ݬ�OǈC-k�P��>��I�޵
�1|�$�lX���@D��%˴�1�F�~��iTU�cƌ鲭�2�HTf�x�a���h)���?��+�)�f��pp��K���>8�����T�R�������K��8`�P�U�eZK[�nŪ5ё�BG������L����"èa1n�H$��E����b��:I��;�r��q1�%*:�
%Xs�@ov�c��Ç ����	;��%u]S3J���`|�l���ya',t�
7�.Q�l=����H�)�%�1}�����3�:�`|��K������+3����
>�r��R��'Z�ۉ��uY���PY���N����ѧWoI�ׯۀW^}��GK{
~����QĒVP����B��{D�K3%�sf�%㿞�5�y��x��W���o46,�";3_�rW�I�17�f�j	�lJ��qz��0��1z�8����ظy+B����ǕC�Y��{�����TT�Que
�N�R8d�8���	T�'�|�CQ�D�.�ӎƵ�^��AO���Oг=lP�6�c���j��&���+m�1�~�]���N�u>>�^{{1���ɘ��|�J�gm裓�'����5t�- ���E�A�)~"�2@;6�j�]�G����Z	���+*7�_�>*,BH�z�3�`y?�6�a������s
\"*D�}�����������&�O�T�ֵ�޶����>�J��O>37v���1��PdUŜ�M��'�C�F[���*�g�e�45Y��c�+��$O�Đپ?IS�*(�k��K��s���t� �١� B��82+b�͎����*V�L����Ũ��IV��a��ݒ$�e���?o8�6�*n�*�)��̙�7�F@�ʉ��!-f置{ͻf��l� h�(<l	�僚�A4Aߕ4�y��ޝ��|�dLY,�lF$H�h��U��,*��}	�h-�ff��ʙ�I�C�3U#���1�+�����ѥ��"�)~X�z��D��{c�}B�d�g�8��8_βiM�N�(ɝ��*86�LltqLg��q�%u�uZ�N<�6>I\�������:��iB��:��&O:}��MP_�[�o�P��4�brp4f�j:�EGg�:�H$�={w��Da�/�<��<��L�N��ǌ\�,���ʵ��#\K�<"�c��$`�<)%�2]]4	��滠C׈�Ɨ�1�5
�� �͔�YK���Er��aM^g�[���\��=����MS+��S�W@Ee�־�,�t�d2���C�z Bd�2Zr�Hu��.���a/�a�XP�9`s{�S~F�$/����Q�BȞ�D�Gi(󉟁�Y��#	�e�����=ۮ�k^�����ٙ����u����"w�A�T�����@��O4D[y�Ђ޸��E¬T���t���ħ��CęY>�`|2J���<�����52p@YǷt�;V���n�=jzk�g��7J�K�*5�_Q�`�#����}��Q������ᗝi�v�DKk�����Y����@�^h���ׯ4[�������L^�7S(�3kμD�Y�YΎSC�S��S��/M
h��%�w�"G&��>Lލ�Y!䮉#� ����Y#���.���𲼌���bB^�mL�pn��/e����<MNɵ�X�f�����bA@�e_����{aԘ�X��yÐt|�G{�x    IDAT9�������/��m��>��I�i4̤ɹ���0��h�T;"Q�9�i��gsK�eI�!��5������+�gI�r2F���f��g1QQ)�R���X��Պ%ཥ���h��:��χ0�:bH�w���{Ü^������B�-�J�Uw5����[�r�p.�˕Ly@F;-�y�rK��"�V��H��A\Fne6
��*F������
���)����\�]x�@\�5�Ď��A���t�<+��w��t�C#"t�q6b��j-6��*��5�}��1�n�!���x���(Wu�J���R�/ߋ�5uehfFQ䕰�b<<r��,Q6�,ax�K�E}�c��Tb��^��҇`�r�ȴ��3m���"�C���r�Է��B��_V�t�%J��N��{�_�-(Į��AJ^�<=U�DNl�D���W�_��@�Eu����H���^*V���I�y�����_����tL�R6�m�͂Խ.�?�84.ݮ}9�Y���ɑ���]���v��j����Q!k�lܴA�-���VA������^����.Ȏ��Q^Z��W�%\OYm"��p*�2�RV=�0�&]N���ޑh�Iڍ��r��O�_� ,�+�I�itG�	+!��%���(�w����ٽ��"�`-���Lb/4�cDg����� �aCt���N�~��k����c��Y�Ǣ�W"��f�V�
}��D/�q�5�wd*����kD^���%k&W���� 5@ʿ�k0�g�y�w�4r"�,:�Z�wI�P�J�|��4vlkf؞�T��dcdʿT��:4n+S3�u�^�́�yD��Y�-��l"U���w%i�kâA��򮰠`a��+�m",|oo�-/ 6L�Kw%e�t4f���ؤ���K=j{ʇ��DW:g�}�T7o�|����tP�qeQ��Œ5>e�L�B�H��g�TL��@b!�@V��i���]L���g],6�����}g��O[�G�r[�
���mE�1����1�${���?u�����	�T�g���	��?�{�ف�����O���hǊ�?Q�
����\�lGP��<e
��Za�1Ʒ/��������OQ�E������R1+���FW\9W|S~l�jyeSi�D�֧-�j���̵�b�='lRU�0\�,��RE��b��F)bn�~�3�Q�Ȣ]��B���^=��K��'�����x�R��lݦ#�=��C�l�5,Cy�S*0X��!Ls^H/	��gs�F�7Jh9�P>���%�� FLe��k����c0�En�P�Gr���4v������
u�q2|��NS�ӜIl�l|B2k8���a��QX�n#�6�Hq@�6M��a!���'�6t��@("6?;\v<쒵`Q�,�Gȵ���3�J�xB�7�h<)'�x�����ҙf@I��tf��`�FJ���\��:��/.ހ8(��4�M:;*�d��$N������Y*���A�V�Y�ҒʣHɶ#1���K!P��ǁ���k�w^� 뜄�~ӓu�*�=�
��eɽ<�ذh�k�;�\���V�Z�b���]9#�6�b�k�����泹�/ύ*�h0��$	y!Gr\[s�K&&I9+{zn�t����l�6!"��8K+.Y(Z���d�&*�g׈T�y��\ϥt{�$םWl�r�]���T(p�(%�|*��$�{�?�h �����<��P99��I
���~�l�*5/�� ;�,}A���d#����
-�;�Z���kA�.�Ŭ����e~"���rt���m�|����d񮑰�'|Jq��^O��"�3)��nWD���?��k��ع��E!D4d�u�)Ƿ$��sa�aY<f^����>P90��G��:�u�r��ߓkU�+����'���F)ݡ�<g�w���&��ǆ��Z��������Fu��ىl&�Ki��z����C�?PD[K��{~"��8d���P���ʘ�y�ɕ�Q��E����**�Y�Rd�ǽ=�E
�#ވ_�����ȭ��[+�'ȁb�󥽵Q-D����Wa�A��7ݠ���A1��C0j�0ݗ�+>��k�$�	N���CFi��oŠ��
�f��Ǟ�;|�\)�l�/��J����������l{����Ƭ�0qϕ�l��y�s딡�̕Xg+�7��P��FE<�ؔ2�����(_�JRk,�aF��T��Zt�����;[�5���5�]�J䋵[��7wރ۶l�f�4�fVm���km�9,���[d	��C�z��%4�'b08�{lòQ���,��1�!��qQGB�B�T�u��Z��9��-�G�"xØ2��ФCT�LWN���q��q�b���6z>�rv�GYeO�kL3���Y��o}f���¦T������v�n�(�46��T�(�pP��)[q�"a��3��e�T�0-4�i�hTW2�D"�DK}��d��f|~�=�A;���N�59%�_L?��tY�Ã��i�
ƹ'�"�ۻ��$��ca=��d�d���y?r���4��~�������I�u^^�x���ޘ�����h3���~LD�B�br�TD:�9j�Xx�Fy���D�@6���Ta�ڵ�3��#�=�9 � ,���W�)��<�P�&�ƹ9?gT�ց���4�!��C��e�;R�'��P�C�q~���g�
8>/�=O��=�J��_|0)�B�.�\�*z�l�Bot��$�C�Fsr7�{�(��j�L�t<N0�]����v9���M�hJ���0��ŠƒC3�d�'9��"FWlh�e����P���L�R�|-�0��b��2?�L�	]���m���{�9c�����CQX�x
/#+s���
��ϐ��|p�aRa�e�����Xx���*S�1��$?�,�6&ban������/�p�{Q�
~ʞi�~�C�|�~��;d{pk��-�"j{�QS�=���l�%wj�ʪj��.��C~�6ׁ�;?�,8�[*�U�H�d&ٚ�oa��$�IwY>Z��A2[;��.�0DÄ����N�ό�:X!�u�����r��Z�QqI��� }*�ba?�v}�ʪ$�s�Ř4a���o��&r�	'���Zk[�l)�(<�!���,�R��;oa�A����CÂ���ǟ|�.�yQ!��f��3^c�iz�7��kMY��T@�V芧�k�q�.�l;��t� �\�Z;�X���F�ź�-8��������c�0"(���.�8�����B%�f��c�7����6&���%���ʂ�C$�Б�F#�	����	9*,d�q�A/K�4c�����#e
�t�^Wj���̦V�D�ґI�,W�V�)���O�7*.2����1U�Cl�FJ�M��5F�4r����K?���w)���jlB�N�\0UՕhnnĎ�ۺ%�5�e��o�^�٫7ҩ,�Z۴`X�o\�VJ���Dmm���M�k����o�HU��)S�s�^lٶUp*�5��M���	m-�R堃&�)L{����5�U_m���{�V���L��])1�:�|6�N"�ϫ�#�\��N��Cc`��zxy�>�t%/�?��B�����o&G<V��R�H_Νyx$H'��zH�,���ߒRvr<t��s����B��;���v���)WTUj\`��E"0Z�3L˥Ս���D�t����ߠ���Y��'�w��pC ���&��?�o���!�p�*Q��\�Lη�;Q�iT���\gŃ����x�(#un��{r��� ����6��Km�.�I�)����G�Hy�Lr���2S���8C��.���\q�����m9�'��&�̯�q$u��U�8	���z<y�=IH���P�BD����$�*�C.U��r0;N|�=	]uy��{.�z�0`���da`N��ѱT��Fd,�Z�u��y?<��$hb!�{,�:�+��x�u`;�H��!C��H��4�מ�9�#��y[[��TÆ��"���6�;jJ{�v�@�;x�ԕ��P<*)��+��ǜ0�|D�8�p~O΁�׃�;����b*"�`zϲ���+ʽ5/�|?���z��+����5��M��P��n�Y�6`�)��	����y)�fN?G>w�y�P]Q��\x�)�Ri�ٽ�F��J�Ǣ��hQCcS��܉�f��5����3��_�6��X˖�;N��lr��r=��\�����W�֧�c����
96����W��2C�$E��
l>k�1Q*Z:������<4R�)6��ʦ2��I�йx �+�������?��6De�W�N������45>�#�sCgu�z�,��\s]�>ɪ3��v��^̸����)�1���eG.� �����QBS*&����$<^�a'r�x,^N8�x�?^�!<.�lܸI���>�a��]W!����֏���y�4����Qy8cƍU�	��ء�_�o���<2����q��1�����J��h���%<��Cػ�̙}.&�?Pq�F2��=�͘�ؓxw�"L<h����İ_��c��ۨ����W]�}%r>�`.���p�'���D8Bs��ȳ$u~�b=<�,�oځP�B���x�	�""��e�]�fL;g�~"z2 ������c�§�ŪMrI��Hc�G�)�	ч���y�M���!/��9�zY:�e�ύ��	���u�zE�u)��<�f�$�uX��$Oh���UI%��eTx�@�U?��.U[.V34���0`�@4\'D4VIu��8���d����q�ü�=p�+�	�,`l
�o�f<�x�
7P"T�b3n~6���eռ�9`��2�J��Y�g�K:3����*�H�+�t�p�����dן��u{�x�!���]Xr���i�O� ��Lʔc< <�M���ބ=U����
P�#պ���1*�!Y$i:�w?���k����UV <6�6
�_P�$�Z���n.�8�������<@"1�7��%�座*���ӥC�#U�E���MGi���d��:e�̨��(��Pf+ �"�^�]��Xx��H���ŻG܏�0C�A�
Q!6fψ�+>�����X|�2,!�S5Ѭ��F3<�<Cm��E��bdwu��TQv�!�����L����F$ �c�����!�"|���?N����h�F2t<@W6��.������������=lF������mM�"��ږx�d�c�vD�1�<_o߁���ট����.���>F��Ni�֩�p/2�}Go�c�����w�*�vɥ�a���z<�F�D9�0u�
>g���7��P_D�&uA�����Ɵ� 21_j��5W̿���P	�]��ć~��BWa����=��|0z�����>���/�@W�6���0!o���m����	-�D<�o_xN<�xA��������cO`�ڵ�Q���"�Q[�"����K�fԗ|�b̜9Sf�n݊?�_~�B�ɓ�ř ��y��F���1p�(5_|����Z�1e�Tq���AcC��ƃ��I��{ｇ7�|g�~2f4^y�%445��e2g�wmڸ�-�ɏo��/���{�F0d�̘9ͩ4����HVV�g�s^~e)���6'�[����&���-@�޵8�س�o��&�ٽ]��S;�/�����P�T���Vf�0��s���r:b�`T�Gp�9����'c���h��-�������-���A}k��Y���:rj1~ IF�A�͔=�Cǒu��X��P�747ĕS��ml���ys|�iGσ����;� ӈ�H�~444�X�%#_<�ϥ�0d�E7�>�kDɬ*C�l�O�7G*N�ݺQ� M�,�U#I�4;8���u�<��n13�rȂ렱��(����^�뽧I�ms���8D5�j%���,p��*>F���s��ѭU�a!;�8��2md�f|?>[|���%��C�������t��#E%��EJ�����w����{��BJ$L�|o�·�����: F�w�t�B��a!�o\�C�3eh�(��e�I�B>Tl��>�+S"�{��
���:T\�)G���?�P�ޓ��3��a9N�k��b��h��A$���h-ӳ��[x�����Sh��ü��f���3	����F�����t�j�c���V�����	#l=/�[�D��|�xϽ��+TT�:k@�����!�9S�A�A�i��K�y�u#>����Z�4��Ϗx�� .��|{�4�y��X��K�;��v4q"�M9\��];�K���D���z}z��X�q�~�}L�2�]y�z�E���;("(�X!Ϧ�/�U��w6�3kt�F�TAi=9O0>���2�5�i���ں��.�^�ˆc�,��+dYX��b�i��M"T%FCHӟ�PD����/+�/�o,T���l=����+�v�o�hgO]�� �\����^46� %v���F�g��\0�V�]d�3�*Ŝٳ1}��hkiՍY��,X�P�*<��o	�RU!�ɂ���c��2t(��}ŕ���#+�]�vɕ�zEtu���͈�rY"��%�X�F���������ضs��e�U8��c��҂E������L�x��|����9g�����l߱��)up�IB,�g���	���ЃE��]��I���;���c��_����i�_q5>_�s�=���-�ק/�ba\vم8`d_��������SO��g�{A�ꚞ�4�̞s6l܉�?	b"�nhQ��kP^^�qù�Uă�A�F!P�`�ǋ�noU���Ν�������(v�5��=���~$��%y��@�Fv^'�by���Ȝ�yB�<�C��w�x�:���Rr`<�O�{R=���Á]�{��/�BC|
M�m�ĎW����S��Be�@�wP�A�:���V2�f̓��x�3@�Ơd;��E� ��$�7g����&d��?�Ӭ�[e0��B������Ͻ��FH9�!,7$g�!�t�t$�"�+�I�8�?�T-��	�O7�OV^T�b�%�`eAXS[+�Kq%�aC.�D5Y��hH�5ƙ`!��ۋ�p�"�ҙc4Z!J�1�H���b<��k ���Œ<�K;$���wp�+g<9w�Y�r�H^ߗ�?7Q	*�"�%DX��c��3K�B��Z�D$x\�+2�B�QZ��(���␤_��l�F��4������"�ҍdHb&)���� �M*���^Qȱ׳���� e�
�$"'��9:62�F0,T�<9�ld̿�#-�q�,B9���>���؈�H�#ͻQ�+��F��0U����[�>� x��ntO6&gV���g��l'>x~rˍhin��w݁�[6�o��"��7H>3)��F4Nw�X� �ϒ��˯VK|�UWa��	������-;$*(P>@����-���+D�k���F3���=϶�m-soR!G��~E��,�s���&��B�sV���)�J���U�(+O ��
/-UR�W�Dѱx���W.���M��)���Ͽk�X�b�	�?p߽�Xr�-7�X_g���hln���:<��S��� ӣ�άH>@\�|���SN��]�{H$�8y��pܱ��9_]�f^�M�>@��F���q�3�Ȫ��eq�z
��/���)פ%���[���~�FuO-ͭ.�ˈ��x�s���`����3p�\Hw�C<Q�P$�4ܝ�w`��/��Ҍ����A����iGM�Q��z7o�c#�,i��n<Dy2�_��'hk�Ãދ�];P�����wf�>������[n�!�x�}���W�NYWCU�UW]���=�ܥ�=y���c�uhn�@YE�k��N\��z��"�44��,�`�T��<����ڔ�3ARm�K�L� Ҿy��p��ߖ��λ��=Mb�sTF3jʠ���m�|�u���TU�O��Gc���b���A��A�=�����v�]]��s����6�:�۵N��LxY�	���"yR����Y��ū��O��M�m����+/�O�����H��	��H�2s��C�!A    IDAT�SH�i��p�DW�=���n���UZ�7�w���ڡ��NQ@b�ǣ!ZĎ��A$��?�%~�㠊�8D�-�U���
A�F�Y~>r��
�B��!y��*�r�`;ZZE��k��w�{ƵEd�E�f�ݹ].�
2�s�D̍H���"��vʆ���,��=TI���ȕE{<��&�����h�K6��=�o�B�������?%�$��r��T��Y!�4I��K��⚒����}��ȸDr+�jD�5?e�t5�����%ERG��[O	Z���в�m�M��5������އk_��Dҡ.�M� �ڢ�!/'?ǀ���5�{�!6�'��x0���g��
����d���̅�9$��\��!Dz��U[�,�XX?�߃�k�7�zKcM�9�R*2cQ��w������u�w�o܏M�֣ԕG������G�6.I>��DD�iLX��'1��98��y������c�&�D���=Q�'v��W�X1b����y�����j��o��^�b�2W�8�/6j6�:u͝��$�r:�F?�Y$�m\�b,��P�F��'�u��?�t��6�����*��n9�����UN�KzVE`�`�%�,����h��s���LS]`Nd0�X���Z&�F�HēhhhQ�-�z� �)m�mv����o�T.R*`xppV��#�4�LhC,��@:�!���>�,��E���x��O�8�|���0|�8�^�6mU��E3n�8TUT��O�bꡓ0j�0cW}��7o�<������fb��;P�؄T6�_}�-F��FC�ӛo��l���]f8�+�{2��8�����?�Yp�u7܌E�����"��b���8��9�2w��N��=�|����`�G�D��k*�n����S߈y����u-mJ�ŒHuf��YYV��v�am��&A6o���S��j����R��I��
��Y$z:O�GX5�wL�C��L��h��{�5Ŕ���`w�к��;�<��ױ���"��J��3Pv	�Nm��!n�Ϝ�ӏ�f���k������|��:�P��	�R����Ã�H	�!D��j� L�x�~&O�.�ֱ���Ơd�<�)#���Ƹ�b�g�0���;�^OC�������Sš�Q/h���3�!i3S��=��D\j�1�H�<l��0�D:(}$�RUU�^=j4rem/+W!Ħ�n��Qcθ6�Pv���r����#kSq�Cҍ~����;���+p�����2dI���4�����!:��)$Kq�U����SZТ�Ԍ�����PS�S�pg�F�D?g����b�
� �#H����C�i��J��AEK+��HVV#F[��6��M�ȦLK���O��<}��#�u�i�����cJB�B��
�f��S��V6�C^���/2�ա$��j�W�d�3�8:��(Uw�8�M,����^�3^d*��6Z�>M��C䵉�a��k.5���}T��D,���׃JPZ]�PjmjF��(�"#��C�a��+.�:ښ�?݃5_�BEY���ɵ�=E2��6�IF�������Ax��/����� qSX�2ۈF�|��d�>�(�]_���������"]_"n!�]���F����ycʽ�vN!�)�XTR�Iy�����ҵe��e��M�R����r᭗�W!*��w6�����Y�zXmM/��q��c��{�-d���,DE��w����l�Mi��лY�U�hhnV�%7yn*ܬ����y�� tO�U7aD���5+eU��<�[� i���i�t�dW���o�h��4����Ze���܂���������6�,�^x�yl��5�Ϝ���;C1�T�����Sϋ���K�l��5��UW �ٌ�}������jjp������sz����� K�,ǣ�>̸��᧝v"Ə���cؐ!8�sq����Ͽ\�`4�`4"��O~�s4�4c�G���Qg� -��IGU{�$����܁dďD4 ���=�{���>� ���FY�d�*u�B^h�l�5���Z�6�.KDFY�5�+T<��wШ�P�b�q�/z����L�i(��c �5n�ܼ<���ё;��0���x�!�_��c���ւL$e������C���u8�$&�B�k:�x�7��o9�l�{b�c��k��2s�T*�b�;�X�ب�r}��kD��S���J��Be�L$��I���8!��i�M��끐>}`t��[�:A�`�O�������>�e$6�?��O�l1�<��:�T�W
�;N�#b!�4qz%���F�Cbt�P�w�
(�v�,Lb#�E]8�@H�Gye�H�$�����@�a�ϵ�P#�#娚����Y���X��W_@�J���֖&��R�f�A�#�y*/K��`��A���P�P���K�}���v���9u�У�Z�B&ǵmJ����u�}��c8��~��PQ�Zlϱm�|�X�ii��`��EO3C:�5������~�hB�����^�c�*���8"��Ut�^ٹ8k�ֈ׍͜��J�7��j��͑V�%ɬ���>5}T|��̫��@����	cp��.C>��+/��-�6��,��/ݩ���q'��W-�y���h1���+"5��Eš��Ps��f�M�#x{ȉw�y͘'*����"��il�����5 ��b��>�"8��#r�`{�D̸O���c��O,�l�Ծ老eW>�˫��
���;�,���u��%!�#��cK{�7μ��#�]p�랼N��,�x���K�d[<`Ef�t٬�Ȍ;��1�5�Lhs{. u�22*o�꒎��io�)�s�F⥤h���?B�H���Ɛ���l٧*4*I6�r'�@.������rRǌ���*>����#����^~+V���-�G��`�C�"����ńq��j%�J'��E�s�Nj}����7�?~t�u�7����ؾ���L>d"�sɅ�����o�F0
�]~9�����x٧�u��(KV���;w��y�gO3|�29���k'��<Kبqv�����P�¨F��.<>w�\����4�A:�9x�pXY�~<�(���^�+m�,���V���?�e�6��G��,��@q�Qg3mu�.�����uw��ͨ�����},�ޘe�6D��x@�(q�vBk\ ��2x���|~�w����I�5ͺH>�/B��D�:%D�	Y�
�����Z��Ӿ;݋��d��A0v	�4��wHs�["	���AqgThGM�!�OWV~ipǂ�j#�$�Q,9H�␇L�60^�b�H�'�I-uOH�sc'������v��$~�1 ����݊�AC��Ğώ��� i��k�i�9��!i$�ڡL����nL��I�;�x�ʴOdk:��m�~�Y����E�KQ��.�k���$�]&(s�g{�%"[��4�H�b4��p�㙕�ZۑI��[�&Dŝ�EL0��P����\���K��#���G<It��8��
��ѨG���<�<T���kOd�B���������!��gh�"pf���̓�#�ܞijr�Z������?����?n$�Mz]..�4��
��\J�����:�
�2��wR1J���C�sD/��!Bܿ��=�^&R�UpF���B"B_�"��ڎ����_��}z(�=���WX;MWƔOT
Rϐ���-I5_
`��z�W���"����k|;�1o|��*�ܸ��U��s���S��+����1�� ��C0�Zo���s�C���({��K)��]�bǢQ�+�|�����DW��v��G{h����(�4�P«R|�6�03��,�1��@�"LĬ�'AӜ}���7�׈�o��ig5N�n�ꈜ]�g��MS>[սqDC!qȬg������_Bȟ�/�a��%�Ö&u�|	�ƎGm��
����v=�U=j0|�p�~�y#��n`ׁn��TWW���ރ��┓O�}�݇U_�ӈ��U��D�&�p����qcF�����+��ر�1zt/���b<��ӂ����y��<�|��Z,\�Aߚ}�6����ŗ��c�9^|y�Q���K�W��<n�������E�b�§�χ��Й��AI?wA�ޝ��hmiDEyU�A�x�Q8�st��N���֖����5)O�s�MNd\�F!��ux%�LY�+̍�̳�lg'�sp2�`��ٙ������$j�<7zO��юW�}��+y��v�Zn�$Ǯk�
v��!|ذ"\���
�)�zx���㌱���*��@I��|'�L�����"s6�b�)�e	��:��\�Mc'�h�@�B��]����(� �f]`@þ��*�K���ڍ��y�t�"Q2,b�yE�d�@{�+^o�Su��� �{�O!���@>�L����(K��ωh���l7QQ-�Φ�6;����%}?YD���/Ho
��P��m<�x���b1l\#s��g�B�
R"S�'tЅ""��P!"�D��wR�b�;����ndc�5n-�^������,
�@M�ވǒ*�Tg�r9e�E_�xER���'ӝ��B��Ұ�a��"��g�4��3e�:W�@�:6GXRf��k,���ٜ%�|��δy�p�g�'C8����v�҅��P�uN�Wt{̈�ڤ�)zo���+T�X�f���e|QIe=������D��D���m�������x�q6c�V�֠�;{Za`�>7&^76�f(�y�/��?��dLA���.TWV��I�^[��P�hS����̺�c�޽�[W�dE�H����y�҇h��91A_��H��.n��~�5]D�D���_�\��&w��
�D0)�B�cJ�烌Kᙿ%��w����Q���>_���0�'�ٮ�F�\�����
����ێx�'��Os1q�(r�&�1����BfI�#���4�{�]�7��QQY&��Mi��-�.נԭ��`8o��F��E5�q֩��L> stXD���,K��:Qv##%�@�����;$F�įI�q�D�4+V���ovKL��Y�f��,�w�}۾�,��C>�g�$D��'���'`��a�ذi�5�A��'���}�޽�˿����+����g�u&F��g�y�?��<*� N�qN=���ՠ���r�<�K>�X�ܤ)��[ߚ����Ěu_��x���qȤqx��w��+o�P���B4Q.b�`�BZ��P[����G��9��H&��oaŊ���yl۶C�7�<t:,���҈�={���^#9j46nَvi������i��Uj<7��&�m,R�0+��B�.C��Ο��<�Ev�D'\��x0�ٔ�;f��3dMD4�����!Õ��G�*8&ї}D����#�J�,�C�Aޮ�����ʷa�A�f6Ӊ��J}/,	��m� ����iCZ���4p�q���aA���T�C8̱��:x(	&$���1m�,.�9�[�[���Q�76�!�h�|T�h��� ��(j��t@�TN^�T�S�/7�}��͘I�����(+�Fz<$��Gk:�"%� A��Y����yT�R�iS�� $@dU�Sy�p3�2�^#"�d���ј*���@�i��1��c0A���2i�=���G��}u-e����vɸ��!f�W��F�|fa��(�{����2e�>K�}��M�կ�H�m����J>^�L	y�k<BD�ʠy�𽥀T����4�l�kyz��zM>�G~�6A|=�Q���dm�'�������7R-9��y��L*�A����δ|	��zR�-�ƭ���F�H�Uy?����x� �o�Pu�/� 6�DI$ޠ�Uد�y?t�'�� ��`!@�B���{+(Ag!ڮ����+95&�C��Tfyo�n6�R�f��5�K�b~<��G�W�y��!el�I�L����$I�:�zT8����6"��׉ąU訮$)?��kknC<�\"еx̠�+��߫�k����-d�]�R|ۺ����g��z��n��i�C��Ϲ��"1�TY]G$	��C�KI����A�Hc�4+�J�>4�b��2qX�{�X%b��ۆ��\��@8�^D2bD�����>�hNG�6�`}���AS�a��5X�r����~��>}��2::[4��ݻ���O?��۷��c���o����6=��l�-�z����O����p����x����R��m���"Ғt7�|446bO�.�5ǝx4�<�P}>,\�8>]��[H�2y���'a�y3@��X�l4�oy���q�$˫F��He�3.I:զ��T�B4��-7�Gq::�ݔFMMmm%4�7�����믾�k8f��q��x�h�o}C6m܂�xHyEǝp"N�>�6l�����b��^Gd<g��e\h4C_]��ksb��Yn8�M�V��b�$�*���L��vm@س,���,8L�6"�K��fJ7݁�w���ZZLQ�qHh�����{��@����E� *���ѰG�%��퍳�:�ƌq���Nk���_�����ڃ떞E��N;�TL�r�������}i�oC����[g�:��+Wk�ȱ�ĉqꩧ�W�^rPmb���o?��V��8��^�y >3*���"7���I'��f��D4��;Ƥ��,���,��8�=Q�܊���╗��bi��18���1l�@u�O>�4>�h)���� "7���+�PI�Ɔ��F�N�࿮�u�%C����yS׫O_�̸fX�1E��P�R�������e��,�գK���F8Ӿ��&�n��e���6���8�kkE8�,�����8����}�,|�)���W<93��+�b�kT��,�|&��Cs6f�X�:��V�@
Ƒ ���+T���lQ��UU�X���/���$� e���E'�V$i�&�J�8��h�w˼����$
�/���s���8@nlJ$Ic����-��$7�0tǐ�*<.[����������^����)��cؤ�e���\�K�x��D�X �)�C�����˛��rv�R_�m�R���@T���!�gT����w�SJ�PQ޲��>r����Yjɢt�'PP��H}4�:x�3��p��F���[
��R�l�-�^}��_�\��7_���k�!єlF�J1
�A~"G��Nn6�^`���ܮgE��N���!\�BE_�Yn��	�9s�e6�H�e�"�c�K>�̷aWVfu:#΁u�V��wfQۯZ�:��q�ɧ���x�����
�^+��8�9t�!�F�XW�k7�Ǧ-��*9pPL�4Q�+KY��;R�$U�|��gX�z&M�$��ƍuXh�O�o�~�w ֮]���F�U�g'���GNAcc�\��,	V -�ATYe����qc�W&F�l߆U�Vi�����C�%?h���,��W�W૕+��k�����F�Ā4�g�΢��)>��֯�捛pȤ���\���r�Y�
��{1r�p�3O=�:֭ۄ��_�����f]n��'��V��6��L�-L��^��6+*�l���a�)ҙ�tm��&+wYq�L���3cW�voT�#��4�RJ��&�I�'�LQ*Jo���e��n���6OA�.T���\��N͓��0���LEaSc���q�q��[�o�6�ݟ������f��nȢ�+�����oĸ1Մ��[���E99�3]8��q�w���=+t���ӊ���'K?�w������0``_�a#�^y�<�̳"X�Ū�������k*sH��}k{�3Nŷf�	�ws/�j�L�|��
q�I=n 6l����'�2z����s���1��J�p���K���hC1��wo��ƽ�g~��7���F/���>��\(��1��ix��W���M�MWV���]��b��Ț����F�%C픍����)����ݧ��8"�Bo3iqT��Ҵc�[H%�9ʷ�ѿOo��g?����Ap�ɧ��#Cumo�u�(��JdS���A%�՜�����{�kd�8�2�&�<#pd�я���rf�!č�fe��JYl/ښ���ϐI�(ކ�    IDAT�⩌�����������zȻ�H�s���D�q����Y�F�Vt���1�3�#����?����\����sG����alB�����&���3/2b��G�4k�~p�����>�2�$�$@�#&�rfT�Y������1��>gZii\�_�w��q[���w��+֜��ԯ;F�9��fP�V��7f�OB|UE5�A����A������~�O�BD�~ˎ��x��_l\��WC}�&n�A�N�e5�&�%,+�O�0:�N���6�҇��2B�;$�e�RmZ��Y�4u��3I�4���Q�(���z��t1k{6m��!��ؑ�;:�7:��sqs<|(�޶-�y�,��~�lݶ%:P��kM�C�mIzCC�f�Ɋ����PnLȕ�y_���`$��d�e��x�֦�@�Z`kӌ����P� ��vTT&Бiլ5�m�g/KT��E�?(Ԝ�,���:��Y������i�T@555��ҳ�!66帎�(�q�6�_0�׬�k����Z]7��F�0�dK}��Wb�՘?�|�s;Ǝ��S�*ch�q�g�߀�X�q�{�a����6�P�9�/�eAJ�24*s���yL�N��%�r���cP�)T�C����g���ש�>�۳��H\k�w���E-U?,�U�JQ��Qo7�2XoS��D躦G����LF��H�5L�nC�+��y�����0q�X��::)u��Ļ�+�Z��+�I'�+�����2Y3}��gxd�\�7���#�� D@����/w�neyf����>�p*�#U;(b�AM4j4�eL�Ʊ�I&c�|��L�o���al�V{h�V�K9��Sw�{Y�y_`�o~��2x��䴽��}��׽�mhT�?݂_����������.�%�\,@�/���7���#��p��HfyP-��|�>�� ��~�5�t���;�j]
��e����V��ɗ1b�8\v��6r4~�o�!$�:��]�1�Fjc��O�����F�92�Kl�Q��8�3-�!���h��1��Vq�1�رcq�m��!��q�?Go�����}��#$f:B��`����F,�F$Ug*"?�c()fI;w:Us�BC37S���w�Kׅ.�]�=���B�8kom�E��s眍K.���������,_���Äz� �AB�	$2��a���y��I�4�����/1��($Cf�H��N�������w|Z������fݼ�QY4�eIZ)X�V�\��1��6����X�28�s2�cPfӸ���P3V���5�I�DX.�*����'"F�-[b��3
�����v�����ƙ
yY��]MS��<��Tؒ�kZ��tm��yEVj��d�%��XF|���F=�f|������H�yM��p[ŕ�}2�Tʚ���3�i)��>$��F=J�&SPC8~�=�d\�<�H0JB��˖��ت�ëoz柿B���J%�w���wt�cǾC�}�|�b9���/!1�D2F�Is���тilnR���sX�3*xYp�P�P[S%ӱ=�w�MO�2�"t����ˏ�@BY4| ������(C�-h��M�{��:e�yz Hz44��PW����AmC,\����d���yȲ���+�1�J���*@�/��e�W@I��.+R5����i�L�]>4'��q�d|"����<��^vF9 ���v+���w,�҆��@"(�Iv~�K(�CU|�����`N� �w�_�݄xē��z�ws����~�W���?"'Wv<X�Qv`�����M7k�~��~�D*�b��I�[Pʨy��W!L��'jK9ww����)uU�&��)����!F�\�����L^���>��mK:�Z��p��ChҮ���K�I���΄���gw�-�������9�}R��7�F�6ri��Q��n4�����cu�Lt�}�]x���x��y`C�hJ;����+��wm}���g_l��=��^>�5�5��]���c�k��q�f<x��p��k.�V^�5=��}q<9�Y���
�;�3@��n��;�K�c�ԛN*i��rb��S����J~�K_]���=��PDʈ1c�c�ɧc��eJ.3r���J��4#��gb�o��p"��:����ea���`~5$JŃ��$|n��녤rT�P>~��an�5�\�ɓ�#��`�s�y�v�,l�Y��>uwT��"$܃zzo��WSS��[p��9z�"�s爫V�{���J�\1>K�C�i����]:��ZZ�߱	Ie2�r�2ZU��g�<�?l���݋C�� e0(^r٪k�zV;����>M�$ULYQ&-_���](Y�P���#/�f@D����؍���:2�j��M!��W�P�'1W���bS� ׊���6��Q;<T����⽴�1�#[��������i�i�]qS�����q���ک�,��7X8v��� "6b'�F/�WT�q�$)�L�l1.y%�[

F�m���D�$T4�S�g R�煅
ӊ) !�&��gF��{k�r"�b>VAv�9����hM��	��4�$�2�U�8[U �13~bf�Q �@!�2���Ő��vH}����u��W�O��7�T*�H�xS"W�O�����5{�Fq%cJT�S�UB!��h�i<��8� 1$���X"�N ��"$���9��wU����:�D2��
�<?�ɔf���?��.'"�u6�=�253|��X��������U�
��@W{���+7���No@]�2]�0�h�����;J5gU�o8 ��tJ�RH�Fu�Q��ɘ.���c1w��E�>d4��aF���,b�d$��/M�Ŭ�C
�P��QB@X��=�6"-�F`2�ry�ߟ@��n�y<�"�î�T���.a�������-����F�6�����y���>w�}/�������I�R���4~rQy��"o8�DYtp��:� �̅g�x�-BN
�QG�d�o%��h��N�=S���޸E��ӱ
�p���B��i�H�1��h���n�í��b�4�V��o�bq�ϳ�cYd亻�B�_~:�oGcm��
�	�g�!q}֮]�p0���>W��[�s�;u�$��n؀�?�F6:��Q����`԰a"��ڳ����u�V=|vn��V̞=]�qu^x�Oxo�:=�BI��<�X`���^J�I<.��{0j�`�}�?�uP=�'^X�<�}n>�L�SΘ�'�~�p�6���;��0n�8�{��hkk�ꁇƇ��)va����8i
Ə��#;ӏ>Z�7�x��
��AK���'�@[s�H��w����זa�1���k0|�p��������?ã��C�UY�Ь�7_�מqک*R,X�����F��ٳ�R�W[[z����.{7nB<���8��s1a�X�+L,��;Z�ZՔ}���X��=�Ϝ�+��R�������Ī�ޗԞ����M��{"8D�/\�"h��qιg�eP����싍x���џJ?("����SC� �z�f�f�׏^�{Ɍ��B��6��To�x;E���a
|�S8C �"ňȫ�F��{%���shy
�y䨊����o���5��,RV� H~��>�7S|Hc��쑌����cfߙ�/�Ī���Xf!�>+_̶��co�"R�Y���ẵ�;Ię��,(0*]��F%G�$5ǵ�d!j�����o)@37N�i5ԾPX(s��b[kp:�J�d��3�����U44h裸�)�,lg��-Kg]?���(���,V��},��{���r���C[oz�_o��?Y�ؿ�oR�J$�غ���-ew�:�yg<��Q]:H�',
�z�Hfua�i��p3�k����䂾�Yt1gf�ae�Y���b	U-LC�C:������N�U9�����H��r�ԇmWO�����I&�>`t�$�A5L����]{�_�l����B�Lg$$$�Eh��H�$`f��h.V�ǥt_.z���$�tl�4��ܰhۊ[
��m�-��ߑ�0ޛcC���(�#uJ3%�i��Xl@�J("�����L��&c�sXcam� 3����l���'��nŖ��ļ��(~"*��:��~�������	:�@C-f�P���~Q��'�Ku��g1�a+�RA�~e�B4�a�<�R����m���p��f0{�;R�Bh2� *Y�bK�Qn<�yG-�͘I���"���D&䨁P���!��:)*��5�[�m�7 ����l@�$�Y��=��6�n�U��.[���t��"j�}�����0ʃ������.L7R��o����a���L����	'��g�!�<�^�]� }ɴe�#QTĈ�uf���'L��{�MN�|?�~o���^r�����?k�D����.�|~?��a��!��x�G�����/��"\���عc֬Y����3g���Wࡇ�ŰQ"Bt�]��y3g��t��?��~�ٳ�]�w�<y�U����{����+1z�X�q���I��N���m��z,���*|�k���a����Zo���iE\�z�/�{�1�"�Љ4��݉}�]z�\;�}=���Sʹ��f���b�ᨪva�����?܏I���3��9�#.؋/.��ٳ�����x���駟��?�Ǝj�3O/Ķ/����}�'N�u7ވ��=r�MR��B�ȵ �Q;kJ�pɬ�� ���X��L���P�i\VM�M�A�E6��\9�9D*��ý��Q�i ��gr���
eٸQ��g��/����s�;DKnn�fپK�2�kP��:��V�d����N"��"����Kid���l>����g��J|6�{�}��$��L����b�p(���:�0뭦:���H�
�$��D(v���uIƒX��=l߹ͽD�h^,z��<5B���v��di���qY3��N��}��oۜ����uC[o_��>��*ݩ��˖��P	~'��E*/����/F��l�(xҹ$������LN�A��ǃ!CK1C7G�Wٴ�}&0��
�t�����@*��	+
�2�4��g]M-r�����X΋�s٤����RŁD&�Hu�z�U��s���9�)+�����tY�@2j�	J��ֿ�4E.�4dg`RnD)؇��h@�OPj}45�f�+4W�t�<��!k�r'>��I2���\|��陦�!َ�s��ŸW��_�²S|�RJ4��#{���M��<��%� �4�C���g���ފO�}��_�m-�RF�ݿo��] w�}�:�����O/�d-���2ë?yKvC��F6�tf�q-�LA��{LF�)w,�6ρ#$��	�3J���P��y����J�)"�Z�7�]�_xĠ��"7>�g�f�Bż0c$fu��^	u_M�5��{7b����������1q�$#����@\���^�իWc˖M�я~�HUT$��?�����	Ƿ�4��C�z(�3���x�}����;Z�J8��<؃�^��˗���"��rR��)}���5NsP��U��(p�I3��p�C$4�N�5a�q�b�������A-`��s�n��#�%�~��>m���W�,Q!��ڂk��#F�aѢ%2O<��q��w���!�������~p3�N��͛7�7��8�3p��7��v޼�$����sq�嗙B%�f�m����D����[�
��y�v�V,�9Nz�w��܊o�^c�5�ƼG��������a��H%�ު՘3g���;Z��d�_|	�����VL�8N���������q���Y|o��x�?���g��W^���Z,[�6���>�l|�����z��g����o�Hl��]x��G%���ob�/aӶmR[R�MK:CP�U��CrD�W8�a��`�觾��*
�t �ϱ�!~٭9ԩ�5eq[)� �s��G����dKa�_�ٷQ�M:S$A��/��le�F�G��lgjS��j��X&oB.�X���[�SvʛJ�j�ia�����0.Β&y�^+��L1B5m�K!�)�r��g���K�z[���M�8�]�	"�nݬ,��ꨔq�� jB4�G<1 �Gff�?yw�ñ樑���؂X"�1ކ��mǗ�Q�{�bY��E�|%˛g�sY�9"b�����^a�A-]����~��O�2���d���E��4]�};�wEi�N(�G0l��\%üO� ��35�aȘ�`�`8����c�f3�B�8���u:�����66���!5˄"���%m���&��Zv���GC��!x����#�ʩ����v�ž���;�WsS>���͟�'�Cs��B�؀S��3d&K+�	�r�nf�B?
&����e��Nߤ��ٴ�T����R|�5fP7c����6�Jbv[09MZ(	+k���g��Ör�$8��,T��r+�#_�[^5d��<h�
Y#�%/�ɰ^7U���]�Kf����菡���'������V���ì�g���ŗ�꒥*I2�ٞ�c")�Un���l�l���d�R[o#�=��Ǝ��18�A1�ܨE�vV��"k�s,`m��#Gk�}V�j�C�Qή��P��я��Ph*�P�y�Ft"�g�����b}�?��>�o��f�}�\��}<��z�M���^!����g?��61>SDTX��c�>�����^nn��G�l����q��������t2�yO>�U�/��?\�<Q"�V����8�u"�J���Q��qcq�nFS}�:�x_����--�L����hljŖ����7�GU8�����3zR�<^}�e,]���:�{��N����+WJ����_ �I���v�m�����_ţ=*[����ǫV�'�������]�;w���O<)�?(Y�뮻Dv�5~��7e@��@v�W_u.��7E�_�b9�=��������L�:|�w����U�\�U�8x�SՆ���o��5&M��\>��| o��6�;�Y8�ӏ�oģ�>�s�;_(?�z�-,\�P�?'�0C�l���Z�~�m��*�s�^|�%�����=r�%7�`�ʚ�G._$j54�S��Bɻ��`��7j�Ji��pT�h�9,���>͹j�d��pz��X��z$p��k0r��3cl��B�$]��,#>cJ<f�d��\�6A���n�|� ���cU��PR6�*%�d���i��Wrek}Z��Q�eH�rյC����Ek�F�d�Jt|�����S'�Oz���Ua�*W	�D�q#���y�PHr�d�Iy��#��d��%:�Mhmo��5b��7�/��y�t�&g�%O����#��6�4I�ǅظ�\|�%�>�ԟ����{���}��)T6%+M����l)pU�p2g`p&�f���?������e ���)q a�j��g�)�����'K�$�a�u;�N� �-�x9#~�����b�w��ʙ�<��U�PHQ_7<N&��׵m��p�٧c��1�����ѯ���!���C�¼V���-��?"7��N�"�Y����}q��Ȏ*�;�PI��B=bm�9����-���P����t��6���D�H����h��0$;͞�&f�7:z�� &�K�TI�ǦL�_�J���Сϑ	���&��B|����1��;v�(�����i���e������uOjjkup����B�X��`!B�y:GL�F��a��P<I�-��
���e�~���ŉ�qٟ�l�Zx�4F�ptc5V���م��^}�3m,�_
m����ų����6�J�ʡ!�"�J���M�з�+��:�O��l߼�==_����*����p�൥K�t�k>|(��^cY��jl�B%�|�2����{�]�IǍ׽߰q�
���{�<�1�[�]��?]n�{�i��ʫ��>?�4\s��C�;kT��O��p0��Lĝ�݆�PPkf���a��U�5k�
֧�~{tb�Fq���~�O?��2�G��1�]�܍Qc�隳�!D���@���ǟ����+.S��Q�&Z�-�u���;��H5v�݃G{��f��    IDAT�#S�X����ZEG7O<��F=$(Sn����;�����|��=<���*T��.�5Z��5���̙3q��Wj]����C�c�!�}�1t�`5i�/|����k�Rq�3�������⦛o2ı��/���=���>�ߓN$�����U8��9:{i@ߦ�6|��/����>!��d�t�����jIi��yJ%P�f�Q�Q�*�5�N���������� �YH,T�sX�8&���C@#d`3Jg��-Gh6crWLe��0�*;���(��?�E]}�W�$Ɩ�8�.^��EGrvu2)����_'8GP����.��T��j�aY�)�l���A/.��b>D�h
G3��<N�:�������B8@_+�&�G.���۱kW��!CG������!#�d�2����,��|N%Q٨߯�����H�V8�E�T{��}{��d1���q�i���y����w=��?��+S�|�]i~���?O�W%r�`��V��l�Tn���$�eQp��grmN����F�o����j��e΍��h�,k"Aԇ<H�u��p��r�G�p��8�Ӌ�j�>���S���$#!7���w&��׉����K�b���z�z���`�����8�C�@��@N�7L�-ʻ���(�璧aF7������G�R���Ee7�J�x؉�������C��r�'��0�_;�H�"hq��f�a��Xذ"�d���b�Q�E��`F��h�^U����)�!cbE�K�,`�Af��.H.L;P�82;�7�V�3ͽ��$�nG{c���t��!ԧ���H@��?�ǎ�;�4�o@��E�|��� �f��Q1�Ӝ[W�� �>	�'�2x�8BRJ6M�y��UL$7d��#T*0���Y�gc,gL��s���y�u6l�F$����9��H��m�HuG�5�Q��C��B�۝�t;EE�����7�s�^,|�Y0�}�E�̳f!��ڿg?��~�׌5w�u!������B�7������_�]{��MD���g߾�J�g�)��-^�%�^��B/]Q9ީ0���i�/$;n�Ģk�ԩ���������;o��y�ŴiSpƬ�X�b���H������>��~��Q>L��#�<"3��}�&��P�����ﾫB�j4�L+a���������!�x����.�+�<�X+d��D��ܢ$v~�����Z�Dro��V]���^<��C��O�8%�&�Eδ)S�~�yo�͛'5�-��@��,��]�Rf��N?W\~�
���.<���8p�?��r���e��l�k:�y�%8����:��g\{�uj�XP������$����}�Ylj���^(���&������>�z�p��Y����GcS�Ȯ
;���bcHn��'�D3�P!�r�P1ϯqR��P�8��F�>̆C��ȓ��A��Ѯ��Bɲ�{��9>��
XГۢ"E����#h39'��4�6�Y{T~�?Bt��%L���Or/_+�ay��˦ qJ*ƙ�z� *�+�6day�����b-V����؜�!	{���x~�s���-��>��'MCc]�t,f�lR`��܌j|��cڇÕW��ۇ`��o�2\U��;��Q��aCP
�OU!��J)f��*��M$����8Љ�g��IS&��'歮�������e
��{ҭ�.��g����'�)��]m�ը	��+W����Ov�POR�<;�8+dOy=&8���C�+�Hx�2�&�CC�/�����#���ػ�24y�l��vbM�������:J��������u���ח�����p������x��V�/9��G� �q��[!�R�4(!���[dZU��<�)�)�^�b,XgB�5g�c.C��k t��8n�2���٠�`�d2-+u"X��#��I�Mf4�1&IT��V�7�-���p�"s�|>���hu)�؉��صg6m܂�{:�FKy��!q�c+f~/l�MP!H�I�6%\.�hoǸQ#	1�҅l:�q��?	�������XS߄\��x"#hr�ظ}�t�zʤ�����Fu��c<�'�9�1?�lg���CW�(J�9~��e�����}�0��tP�C��J%�_���4M���I�O�E2E�:;)(,3+P�*1�>�{�ضe�xm�PƩӏ��7ߌ����Ʊf�j�Q���՘��;oC=Y�|��A��9�nomƝ?��F��lq��;�������5�V(��+���)O�T�H��������$Oe�U��I�%��#D�*�B�"C'F��o�G�܍��j��^y�U��i}mK{���G�{�y=v��,���N#��#ZA��eW\��/����>߄?=���k]��]u����T���&�@~���J]�:�lf�|s���3�"��c` .G����u�Z�<�~&�g���<�K/��6������{!@�^{-�M?A��/��%���SN9�~��zw��ٱ{��.�1B�q���Ux	�馛p������oѢE�u֙���\��٩�)Q���^�lð�A���`���{�\<D����~�����<eΜs.b�,���&v�萚�V�����2p�Q�|��֩���p/�%���+�£���j��e�f�yv�/)��Ъtl�(�dpT�E<c��3��k�JN4Լ������o�!!Gu#��0�c��i�+�c9�'���l6)��+¿S���e"�b܎�-�_�g��Da6�(�ܰxz��35w�8~�����{tyX�0Fa�ؑh����Q~.�T2f�XSa�V�ĸ���~�9��Uw=��*,~�U|�y�d�􆩫�ư����w!�A������P}K\� >߼�lٌ�a��1x���E������O�}e
�m�J��{_"��N���)m,bĈv�8i4jB���۟¢�W`��^����i.�q�����w���> yͻ��A$��oT70�r�vL�0
9�r��>�C�3��Ҏ��/6a���H�Dªp��Qcn���������.<�L�z�X����'ѱ�+�_��Pt�O�T!S0!m$Sᠰʷ�R\(�IR�d84G�`4x�l�Is #���3��g��DT�0���MV#!n"�������h��Jh1���Huz�wq��8}
hi�	c�se�������"���~�7��;���ql۵_n�)�>n��!��~�e�mи��8q�<�T�<.���j����@�خs���	e�-�Pv���E��W�͕P��
O(�wV��_V��ڱ͖l���"*�,c$}����f�6�#е�Y4�c���w�>��H�BCC*$�I��M��X��f��2��-[T(�e�p�k,��f�ڋ�q��w`˦�X��B�,&/��R)\�����������ln�_��>��X��G�|��UJ���wh��2�ں}�����אہ��g͞m|}P��zk׭� �Ψk.�4��+s͋IR���!�QÆ�w݉�pDʫ�֯�s�-���I:��;�\r	�u�?�Q�ſ��hԈX�O<�V�X-��dښ�Z�����kK�f�jT�ֈS�������7O��{���!�,90Dh�H8�2e�����=�x|���"׌E�w��㏛ X��� ����=���|�;=z>X�Z��jtnjiÞ�����g�m��~X����B�{wn��nL�0N���|]l4���:�yx8���+X�p!�M�&�JCc@\ظi��*���l�}r,�؍+���+W(T�7ޤ�˲�����W��߉�S� �72���.�U�^��&_"�|�y�{]
\��W�:�dШ��yy|�<DI�%'� �xM����c9�R_�E������m>�V@�='ZaȲ&���{�;��#�S�9p�):��Q�+�`����%ߟ2��}n!ng�LJ�k�:�/������1eE��o��H���xo/8<�7p�)[�fl�.�{��)�c�}�B*�&���'��6�X�a�t!�N���V��D���!�~�	��X��x����+4x���X�z�
66��5�7h�o@]$�R>�J6�Y����,9D���mm��d���/P�҆!#�����~�����+T�Z��g���T��:��("�w�������%rع/����ys��]��_u���KN��zpy3� V=;�	S'�QE�RU���o )_���^��������;Lv�TQ�P�%P���&�֖L�0��59z4��<�?<8)����荥3υ-��e�m/j!R��8.�����P��2���P3��H��t�@5��*��gE����!r:�D&�H�u����x�dmӛ�P@42�C���?�F4Z�TP[[���z��矼v0$���>x}ż/�PCc��h�u@I���������[.�ȝ�T*
H�p�Y�9+X�zz:���Os��:��ڈ��:+�g�X�9���mF,]���1��ax}�}��T�X��b]n�<pH���M�����)L	b%�ɞ�"���H���fCӂ��)2����>DEG>��0C���C��kbj��X���g
);Z�k|���{>n��v�p�� ���O<i���*lٲ�?��4��3N��_+�����g�7��m-���7`РF��:�ε�t��nq�gh\ϟ�襗�ʒ��E���Z�O���:&���p�N=�|�JFl:��+�����nA�C��@�С:l^{ml&O��[��=Ԡ����0��M��kp�)�"��(�AM�!���|�u��u�,\~��hh�����*˖/_�u��I%E�,_�3�T��3n,����jlX�.Y�D����#�2�W�HΙs����˗k�{��s�j��o����q�E�����n!D�lV���A*]�-[���~C��n���M��ܯ'�zR����c���6r��l&�g�����?C����U���g�>:J?+��܋�6}_��^P�CߢL���q�%_��a��7i����0)3E��H���g�5�A!+�#��k�Du��-��G�%���c�b,�i��N��0�1&�i%K%i���Z+��G*�|�{��Q���,2p��ظT�0���VȢT�R{���<��`P�HȊvaӃ�P|"�@@�Lg���%�<�6�>]{*�h�GD%��K�k]�8e.����9Kxs���q�Sq)��|Q���4��8IH�s�^P�ˌSf"����W���`D"*#���!�5��Z���}=�&��K8$���&0����6 ZۀQ��≧���w�9�w?[��AT��*-Ͻ�����t�����NW �Y��^�(�+{�̘�!t~PO�����<��0��.��J��w���'+��yT<��Sػ�S������C��<�V�В@$X�XЃZ��P[D�YB�!A~����eW`�	��_=���j�πN�TQkn(\(�5�7Z>T)�����A���p9#�̿��\����UႵf�B`x�z�����x\��nT�Y/��8ƍ�Z*�n�VU���hIU�ǉH؍\>m�dyO�.�]�N����	��hD�� ��^<�9�!�g�~��w@\#��Y��0�T)��hW}�b޻o-]��ׁ��0�!D�~4���O��vC@�\&���Q���ص�w���p�߇#���~F���q8�nl���Ќ^��+G$�v� �9G�,�m9$�y��Je���VAƃ,���d*�BAdXQ��f�,L�.ZfR�'��3�i8l�"�0}�:v~���,b9={�d�$�q�G�̙�c���G��ׯ]��?�B��O�������Î��꿎V6mڤ���Yg�R�@�����;��7He)�bZF3����!|�,ƍ���<K*�\*��hD�)��E�4i���h�pw���G�5k&�;F�[n�{���;o��;b��?�8�,2X �Y��}�):�׫����?Ŕ)�QˑE.'e�>|��w��1�1c�~tʃiz7�9l8��1Y����v4ν�^�D��ČNĜ�g����)���ӫ��<��=b�qo-��ɧ�l��Wƃ�E�'�|$��g�&�k"g���l�5Rva��)�6�쎑��~�7n�J�����M��j"^�|�s��)&M�)��������Zlܴ�u��E�%2��R.g����q���N�if	1��
�s���6���P�x|�	F6\=�-ʚa����h�C^�%8b�v�x�.T�:h�F�P����*�!scy/����@�[��co"Ύ|�rN�%���.�(	��5+f���kLB����=���2�{Y8p�5��v��/~�'�bq��7�q��p�p�ɧ�O�x�b�$C775�P�{�y����~��ShO�
K�h2�N<^9v�^x�}�'�6K�嗗,��]He3`�n{s��w���c4e��=p��3��>��@���5��knǗ{�;n�d<�伵^����
*�J�3/��e<�v��	$���,P��;�4+'E1S(f�m��%�%��W�r�(� g�	!e&l����u��ڏt&����
�����{@�J��p��%�3I��ƹ���=��M8��ؽs�`��s�)�O�>�/w����e������?��.��E���iP��i���U�p�a�E@�B.L�E87�7G�\�^gg	���x\�g'F���%�l��x��wEC Kʱ�FQxnڅ���7���5�\vqF��C:�SǮ�V>�X"��朅��G'`��)^G��=�����5�1~hڪ3�E��$]S�ǟ�05x0�)�?YD�Bgo
ݱ,�������pC,Z,3>v��Hj"�֎Wg�r-9�P�L؄�Xj^�c]v_<(�-*��T��K��fAu9*,(�Qag���
Q3�F�`#3��Fox��2�~HE�u!����V2fa��y�(���*<�����f��B�w3�B~	.���+5P$`��̬����,I}��pN�^"\����h���!�O�����^l,L�J���'\N,^�������po��,�O���"��E�q�5�I�Pf2r�6�[c^n�<�y�A��C�!�R˹gQ�v�����[V�a�qJR,�qX�����y��p9�	���Ktu���8j��_'G��8Re�ϵNgZv�|�\7�"S$"z `�2PѺ����R��GmC���x|�36�١Ah��b�ϭP�.�)I/Ɉ��	rL
�wqzX����˧F�ذ�u��\#�S�Y^��^����(��@�b�Hn�7R�iu_���CQ%$ӓ�F��$�o�0���"^��H�9�ZX(�����0E����^����<�yX�Q iN�A�Rp�L���Ȍ����D�m���7cKx��pKF0pP��)�k�!Z�3w�$�)Q�)0�T�-�r���O��iS�c��Ef�^��;#����:�L(�ty�}�'�3���m�8y��*�^x����k8�ks��╥o`��zV�9�
���6�!�v����\Rk�g��Kww��`��1��Ջڦ&L;a:�=���J1}��?�����+Y���w�5^�_�wF�,T�pS��MV�c��N#S�kQ����,7��j��F�TPv�t�����dR��Sp��c��q"�-{������j�hڑD�cwļ ��n��dv�PS������Tu7
��vi��{�AT\&C�K���CP��Q<�� S�]���p#bמ����GI�ƪYh	fb#ډ��ԁf��Jςڶ�&r�1fɣȥ��:���P����H`��8��3ԱH=�p#��7!�r������]mr�/J�($��۸y�f����7B�'B�
85���d���_�~J�P��Ϟ���=س��mo���5�Qվ��ް��p�;�D���TW��2�8�}�7�dԷ��/-�K�m	^�֫NP��3�G�i  �W    IDATư��Iζ��,r�A6��_��2}o̵�=�f>d�ptuuiC��!�'{m+/ɨ�X�Xd^A����<�x�ҟ������3�h�D�B�?	��I{|�h32�4�[�N���6��Sk*�+03��A�h�4�K0+�d��ԛ!!�[��١S�ȭ�[q(L�.hT��#o=�F���|��-dupR5��S�JI7C���m4Dt@)@"3|����w`�p+x8UWժpaC �B���ѡ���*��Y$��QDrMع��|�����d6���:�1hJɎ�k��~����G:M���?�54�#����f�k��T{�)'Q.y�H�^����vF#H�f��Jh��(:*J%�x���]?ݻi��F�t�i��`Hn�q�E�����{E�`*C��S3ɽ�(�l�H�P��Jp����4�d�_6�"�D�Y]X{ޑ�r�@к�2v�zP��dUʁɏ���Kᢊ� ��ڋ�?��RrY���k<�C!������	���l!�T��h>r3�3f�K]�fWE�������i��؍����͐��7����U��0 ���g��S����P�F��#d�IeխLK����G_Y�G8��3P��k�V��??�9s.Dc�`,~y	6lڪ�OK���f�� &����#��!��WEM],�Bw�CGb��	ضg��Z�`�z��u�B���՚���������B��D�a���/�.�9¡LɅ"����)>���t*�Ni��M�����TMTJ��#��i�@�ef�0�ĥ�K��G]C�:}���p���],VRY�.��n�o� )@ֿ2��Y�\G�9��bW3D��u����D�g��w�\Vv)�Ȅ�%��6wB�rpd�lLrQ��=�U�!ٜ�!*���-��_���fj�f�rt� +rm�T+�	4Ԇ�K%�9�	��e.�::0n�H\p�y����m�
�R	������ʑ��U��l��{Y�0+bϞ=r�l����^�îC�<7LvR�w���9����3���.ԅ|�9}2���aTk�h��Q��G]oʒӅ
�2�=�ߟ�ޞŲ*V�M<C�`�����F��A�f�.y�Z��Gx"|2�ʒE2��&�ڎ���Jɢ��)��5��P�����*WX�T8*ٔ	�&�IhYT��δG��c�}2X2�����1b�0�|������Ĺ70C�3'�yJ��Sz�v��O�P�ۧ���X#�s.[BO�$�\K�QἼ�Z>7|O{�0!�L{�]tY|[���y�$�f*y��H����ǅZ���C�9�?� 3<��]�"�hp��e������eI�����X(��B6����d��і�a�Q-n��I����߯{˟ǵ���6d4낯�4r�L$U�s��f�H����w��Pc�C��P�<"uVn}�AJX���'*���2������ef�D�I�X��.<0�f�h��������RA:��*�둡���/h�U8�#*�$�<���Vטh
�e�y"1�F^$lp��(����T��p N7q�r�!�����KD�_�,�NY#��H���L�P�7��(*�{���Ջbo��EoAymT��X�F�Od�?�cY�(s�̘�/�r+��ҧ�|-c1��X�r����"G�AMM"����H�2x�8 �0�#A��iS!�2	�~�
\n?��p�7/����?�A6�Ѱ�؀��~"Ta:hmm��>��M�D&�%�����>��_���'��'��ǟl8��]�eP2�>�'x��q2�,(()�Ʋ/&���f�_U�u�n@0Z��3�c���+�_}����?��7)Tv'�M���U��t �
�JN��8]�к���̛�]e�}�1-6n6�|�Q�/�f�$H�K�X��Vt:���P.��� &B�t�e�"ک8�ƌ�����<S�V�-�%?�ȥ*�\K�K������V5Lx:>�N(��ա�pFJ8�iP���!~܈	iWd�ύ�d
r*ȷ�6&n�\�|�	�r3�S�+ev�D�~�Q����#�F]UX"�|�t;�m!l��q8夓1r�p-Fj\��y�Ox���i&]b�hl���4�b����E%׉lRtB����,(�8U4*��R^g	MUaL=g5~Z�]�q%Q��� ��!�6>�#i���GЗ)�/tN�3Qġd[wu�e�DD�G��wV���D	$����R]�T_�J`�f�!�hJ(�3ڜ�^�<�9��դ�RF](eEqd|ßI��M�T���A��(=�EKq
�bg�h��P3�J���F��س�u��tk��p���#�* �ɱp"	�\J�y8�8Hǳ��)�Ac}T�{���>>o��`&�z"�b~�œ&^��T��2 ���)�:X��|>��Ϛk�d6���];y�<�|F���;3J5�+F�şæ"�4�m\�+Q��� �4�7YJ���<o��i:}~��U����Y�D!�~!?<���k�<S��nGQ#��뷷o@�	��D�|>�f�� B2M��.�����a��ȼ��s5�M�`�;"RZ{���yd6�G���PU�)���.?�ټ�*.���%}wX������PrTj����^̤gU�󵓼�}�t��V�}*�sM$�hl��Lr@��0�Pʣ�q�a��q鹠;5E�������ا䀣Hj�񒑧����|n�,R��W�U|)�����s=�;��А��/"!�Dc��`L<nN>�T464�±R*�Թ�=���{�b��]ؽs�
�}~�#N�Z�`���p�i���>o��6z�zedʆ�����*4�T!"�b�$�wT^R�>f�h���|�=��f�R��%�c¤�x~�KX��gz���Y��rg"IB�B
$�:�����}8�u���M�1q�tL=~
^y��u�R��ŏ�r��x�rT���ޗN������#p�+XJ�"=1_���_U{"�
����4�ea��N��Fo5�0��65"�,煆L�LK"�0�
��݇�+�d�D� �_�P>�]���ɥepSf�S8(�P�'v�^3ޠtS��7��d�����Ac�~�H�z+��όOX̰P��F�u�Q�a������lS���dQ���+�aqT��Sʡ�YBM���.i��?�;���,cڤ	:�M��Yg���p��6�B�ȁ}��w}�B�XHvuwc���� �L��^�tN���&,fb��`=#�I��!O��T�!/�����*�T�/'Q̡69{uᩘ >ȄЉ�8�K�+]��X�;��ɖT����z0>�l�:��]^Tӻ�
&��}�Cq.�೑��̓����D	!��9��a��L,,�s�hk�lcԪp�A���|%�`�&��8djx��2?��G����� c7�Ε��Q�	r�|*���"=V���dA�<�Y��3�q����`U���\��B!*�xL�
>�,����;�EI��ק�'��j|M��\ޒ��g�@��r��s����*�T8/��`��-�ʠ#dSI�l��C�O-sD3f5P<Q~�|I���n���Ȍ��r�v��i�޳-�B�T�x(#�:�T�Ҧ��H W�����A�rj��ؘ�����h�x�o	���l��8��_8z|�{���s\Fz_!��a<��zd�Hsk���b)�]�U��O�FU�X�� ga���Y��\�e��v.�R�R�z'�!�$g���$0W��Tڐ_y?�+�rd�}�;�����O"DYʄ�i�D����ߖ���B�#!����hǊY1�'=M�o!�ZF]m�[���˃��&tw�Ŷ-_1e�B��N���Ju��G����!2d�L�ؤ���(VWw��Z�����	�����#��G}�g�^*��J��s�ۋ��#��>�]/�s�7r�������J{}_�/���>q�D�8��ڋ��XGمH��!���wW`�ǟ����Q_EC]�$���r�\�P�@X�!�܃�	̽�7i"^~i�(%�y����:���J�~���O�����n�\��-۱a����sdr@&�D,arFx@j3�:��nD�����
ͺ	i�O�UXp@I�7�A<5 ��t"�h��M��W�y�E�.mR�R�x�8=������u��Q�&ˍ�_�L�5Ӧ-=��R�̔u�S�ˢ��I�~��WǛH���P��H%5���C�
$����6�$���50p�Dc�T� Q]~�2�;�oƁ=;�<�>w���5���O�8AŅ��t���Ԙ��)h��H"��z�g�c���D�d�AX��W���l�G"3I�܆x��J�Z�Q���z�nm@m���:PF�[F�瑷
�u�>�%�.+`��q��D�@�
�q(����G�iJ�A��qP\'v(4��׫Xa82�-����T���p�2�����b8������s���*LgB抱����732�RiTx���v�X���� �"O���r�<�������!o���(˄�8x�Q�J�?���h��r������\�Kb�a��=��g^���2��~����kIϯ��Y_����;J4Vq+��6�3����˯��:Ό3m��g��`��25e��m��)sd��cP ^'�&K.n�[;��~�6W�j:si�2�����9��S�b�ϴ6��Xcb��-��`�{n���ٲ��y���#
��#�6���������I�E��X��x���x*�I��D�*�K�'Qb��#ϡ��9�ܷ���	:e�#.�9)�(_�m�B%�"���_A9o�g��m�yN�4��v�߇P7�Gf�����YzI!C^o@�YUȇx���S�h&�F�4w�@&�"�����1#���GBUܸ�#�N���?E��C�gSȤi�QFӠF:\^<�
q���jTxhϓmY� D��>���B��W��F
6�qɺ��ǘ�V7ԉl�����6qCvv�����+WW�q'ߋ|&"��&�	��:���.�A]�˿u���._�;;�r�Y�IA(�C8���͡�&�f�Ea��]e�/�A,�GN�>{�N��%�.�����ůR��T���g���ʷ��� }-�kk��x�ц���s$�$$l[B<�����q�����h7_(iVH���o�W�%>�� ��<^����w�q����@�-�V²^u�\�5a��{{c��BQ!'�xWD2�GB7���*$�{cҞs��`���O�mV�TIm�����v&���*!�b��iI�#�G�(�J d��Ao<����-��w�pd.
p�?�	'N��ߖ!��Q�D�
�o\�u̙=�uQU%�~܄x�p�gq��@����cߞ�x≧�삅�.�n��'�̈~�H�U����lq��x��i�Jp�r���U�T���A�<���p:y�z�Ö�Z:�r�9Лʣ3^��C)�ݴΪ!pF[�Ŏ}BpYؐ��Q�C��p>+D;(�|�{v~����(d�:�ص���*�*6X�ڇ#I��P3Ϡ|R����FHt�㹢B�:�ȏ��B��J��t	1�l@6�p��)�-[o�XЯ�
#z4��}��%\�0sD��
N�|�H��'�������mN2�#�A,wu�m���ZFv�(�>�Y��cBG=j��0���BE**��:2^:��DD����1�E�����@G��&B�τ��H�7�]�2\�^�@�k��q��Yd,ʙ.���u+DlUq�l�d�p�k�o�E,��#��ۯ��N��e��r����[A*����d�}�#�~<V��.���k�HU^���Hf�w�G����9s���2���T7DWX����%��2�\䬩��	��*Tx8��8����Tjr���Q�$���>�BQ6���B������j8}A�R�q"@����ΙTn�_6�y&(��#7��B�mF�͆��%4l��V��={�e���ŧH$dPx��;z�Q�+2	���7	�>+��q#�� M� ݫJ��lB2W����L�N(FMC#��
Ǝ�(d��N>JF��TF��Q�S\$�;2� <{Xl�}z�-����s�Ek�`�X�>�nۮ@^�Q!����yc,�0N�Lɮo�Qc���{�it<�'��gL��o��a>�s�+��3��H���_��'�����f�N�Z��3��`/��+0�,#�&�8�D��J������Ĝ�q?����40����Y$��Q��`�f)
	�=i��T�7~Z���C���_fc��&ށ�ڨ�^\�{:����7������Xl��� �N�HE�:�
�L�ر�
Q#7�pݐ!2�"�$.Au��:�!t�ư��!l�r�`dV�T��>�ƍQ��J�/����`wL.���W>	��B�� J�~L3�Ϙ��K^R�f$����s���.85��n8���O�]��ȭ�M�Gv�V6�Ӊ�;;��Ï��W_��:|��,Z˚�Rv7^ҽ㿑8LtL]��	!� �h�	��>�j��a7�j���x I���j3�e�Gê|1��p�@���4��P�o܃���h>��Kc&�h�u���;��@J��ItT��ڌo_q��<���؍(ɚ�T��MvG|��H2�	�d�h�#$RE/LAa>w$k�B$l����9K��[ʯc}T�=���BEEI�Vx�)L�oˢɃ�ݸ�p� ���S�kv�^C�>Q���co�ɬ�<�%��~�7�"8��05�рG!��	���Gr�)��PX��Rᘂ�~�,�͘�# C����D�d�d�UCD�"�Jv)��p�����U>�XŇ���?��
9����3ƃPM��"�J�uԴФ	��m�G4�}���%K6o*�j;ܼ�=�oq��T
m�� � �IK�<�ԙ�O�Ŗ/�^�n8�c��QM�<!)	�P�UD�����9e�iJvR9*�,��E�F~Y:��Q�&�,�t�X��D��2�$͑���D>M�
`�����B���"�^���3)��6�+�I�%q'r��� �,
����sDga����`�>BmMT�=�Ŧ���s��b���hok�N26�#����}R���
1a�|�0>��=B�ww!���}˗��m!	w؈�����x
�tvb��L=�D�:k6|v}�C����{{��`S�̱ZCc��JfC}�ɧ��}�s��76a�{k��"�Ҥ��_�F�4�.W�L����ʘ����H5b���؋=���Oôi��w^_����ǥ��b�[�����oB��ܝj~���Lg
W���7�@4��sf��ï.[�}�̖�˔5n���r���P����u��.���M�5D&����#��N8���?1�Ɍ�g�|7}�a��p�i'���N�_]�C<	|��X���:��M?��֥�{`�H��7J{,�PX��<��|9Ur"��+���@3����r�9f�6�P�$3F���KK�z�*1�i�s�磹ك�^#�s���Vn�cO?�8�<sزN%�{qx���cҘa�2t�3hi�Ž�ޮ"���6v�'M�4wv�:7^]fs�>v�,y��޽������L �ќ�s��ȡbH[�\�P�[g��*�c�U��QDku ��!*��<�9�RE����578�-���"]�!�%�։��,�nއD%����]�����fV��ٻS��V��@L���|�v�٧��`���U�A~C&G"�� r��?`yY��AUx�Z��G�"GL�_b�t��@�3Њ�����;�ݧ�23gzW�]�lٖ�\qn@�� !�y���<���r���psoZL ���r�%ے%˖�{��>szo/{ϑV���z�Z^n��̯|���?����ݘI��f^[ꄃ9i�dX�P����	xͦn�o�=� �b��LF�˿�4Q$9�0��D�k�ӉT����|e�'��D�?��ׁ�ٔk��P���ڵ��X^�>`.j�?H6�[o�&Ǒ��h��    IDAT}j�X�Z1e��p�`�.R��t�`��1���G���\�b#~�FApd��1�]�0�
�f�|r�Բ�j���a�:�� ��N�����.�lµg�0��06|/��a�C]ddC<^?��>\���C�tpxf��0�d,;di�P�)�A81�]p��($�i��Udw�@�z��Q�=<pQ���/��82s�($g���B1;���fp�mt(�`��VZw)�����Zmu�K�V`�݅�ÅL���br6�jT���v6lX�eK����cbTh�_�p��[s�*����Њ��A��R���ۍt*�g+�6��p�I�?$ �l��I	Tda�ӮYZ�y������>��pݖ��_�,�'f��K�ѿ`1��:�H[;/]&Qx"��j��2Ç���n2%�Y�77;�χ����F?����X6���4Sw�0MN)xP��a���{�E�V��d,�Cߖ�nªK��K���%&�����d�/����/��OV��{~緋e�#�l������݀�D�w���Z���E�*�L8Tb��+�}��Fι�Ad,��;�<Ys�H�j�l�^'���[��ߺC�cػk�����
��掝�=�ށ[oـc�Nb�h7�-����O?�2v��&6^}5>��u�N�S2%?/�7nي����_�._8����s�?�	�=;(���裟D�P�ηޔ������$��O<��g����k�hkQt����
K��_����mێ�d+����T����CQ���
�4>�m��]����n��A��fa���Q�cC�����O�$���B޸"��?��}��p��b�bH�k��r�X�s��v�D�~$X�[�U�t�%���=�A�^DOK��A�~�q�e��}��b�8�e���l����1�f���p����^!܄�EKKe18:&:T�CtrE�����fvl�l�͍QK!��avr�#CW@㰥(��E��6��}�^m��G?��\wk�ى:e4l�%Ƭ���6������=���?��xpswM4x-4��Xn��j���@�8�j�?�{�{%�_(b��D����є��y����AGR}lR_Rj�E��Z~M][Q�V
����7m���� TcR����U�#-\ш9��!��L@�0F�� �6
���� �RC}�$�����X� �e��zoj���P�Zs�������~�٨Y�?�o��T����*W�]�9�`Ե)�Y�.��%�v��6H�3?�!ddy��~�>?���9u��U�N�Bݠ4*B����d��E�#����oƪe�M%015�k͵�����A$���f��#�*�YJ�ʀ�������H���	�]*F4[��q6�A"_E����tN,K�jC�bS�H�d�p�:��Ip��I��n�i�c.\������7�|�2Ѽ������TN�>��"��q����=�j��'���lB+9��V�L���~;q
�,��z�t;�أ.��������<���.�)V���QL��C9�c5�d�'�p�NFQ4F�ށ8r���8<F�U"��e��c��9<�8�H�3:2t1S(#�"E�F�W_sV�Y���}r�-���m���_Fe8^m|�ŝ���?��-�X�v�!'��?�㧇�/��F;eQ'W�1{���p�l
��R剗M�8���Xb�r�����"�2nܼ�]ۉ]o��g~���p ���k����3�}X���?(++��%K����������O}
����SOapxDu�|`�n���s3���3xs�v��Ȧ�[��>�<Ο?��nߊk�]��{���^C4�քm�[n܌��i����r�9��O���"S�jcv�"�(�rh�M�������J��߃�츔��b��݈�~�x�V�4"]��u�ᕎ*���L
�{}>̍��IQE_6|�o�������bq���
�rM�e(v2(�s�Q�����
�ث)t�\U���-EtF��nm�؇?uJT�35�:#�����f��)�'�8|~c���^LDS�7mN7� �/Z*1���4ZZ�1:1��gΪخ����~+^!]z�}��8�$(j�c@<uqlB�f
0��ր��R;!�7�z餲<k�����~*7vٲ����B����I]Dk�ʆI�&�*ʚ��T���Ϩ砘^��'FT�s���r��z���P�N]��#<��? [��"6�،r����{��kd!&ƈg�_���Ĥ��Fk�ꮢz�K��"�-���dS���Z:��=\��#׀��rʊq�|�UW@�0�,�������W`Ԙ]A�2����q`-��3͎qܒ�Vs���>����P�]�Jaf�R<�ϑ0�֣S�2�װ7�+E�lQZtKK+��y7N�ġ�uzvz�
'c��k�p�-����󷴴���1�)��¯!>;�緽���A�P���m�Z�*����	`Yw3���h��U��qm`9+�z��Ite�w�(���l"���X���DӪИ�+ZPu�����-X�����܅�8z섘G�LO#6;#����p�,^�X�B^�	�K%�051��Ft��(9�,��(Хɀ�G^fEQ��1f�'�9灛��|�+���Qv��P�z{/b�V�]��o�	G�����$�/\�#�N���x�̺�;���A1 �>i@%S�L�1<:"���M7݄��y5���g����ON�[D�����eZ�9�`�c &�W���YLL�(����6�՗�=`�d������:+����¨\HV[�m���d&�pCKCxޢ5�pqp���\��F3�i�T�q�q��)���h��vQ�P�u�>y
#V3�_���������}���5@9���$&�&1pi�/���KX�b~��,䝌�ѕl�9�~:|����������7����˓Qj0�T�|�J<��ð����?�6\.����ge���G?�����<�ښ�OO����wŲy�-7㓟�8^�-���k����nז399��/���8�9t��s�!թŲR�>�O~Ak	��z3#��>����?�y��Q�sΛ�����:mNgO����^�%�X2�?�˭�Bo�(��/�dS�򛿅#��K��O�TZ�<2���	0�����rl�ʥDF��gC�iAG؇[�}��h
�� ���JȜ��nNx:[�t8~y#�l�n���_�pSD�v�_@e&���z�SgϨ�n^_��nl{�E\:wScð[)#���RA��.�Q(:��Y�
�Ź2&�m ���M�f�'ښ�ń�} ���fO�@vÜ���brl��ư1t�1ņ�]�+�U��i�� 6n�5�Q�.��K�DZQ��zژyb���%��h[�a~m����4NWFu�R�!Tۀ��&�8�2�+ �
��=�ɫ��T>�ISd�g��E�\{�(b��G�hl�\Gu�j>2U%�V�A m�СRwa���!��ϋ��1��W�IL]��7B��/0ck����#���f�3̗y'� �׏�M�Ђ+q�U�?���ח^�S�� ���՘��]��N���c�Tܾ��YH�s�`GEzk���ni���B���Ɗ�nL�����:y}.�214��X9�������|����a e�D�[���g���لN֦�x��t��$ Y� Y �����a6W�\ނ�dI�V�p���x�fL��p��Y�^�m--��Awnrm-mX�bŕ����iIX�273���n���K�>z�zGפ�. G{2�7��ܿ(X��zv3Ԧ��ғ0v�L��	��&�p��Y�D��e�mZ?=���>���	zݍ[�N���e `�|"�;���׋�y�c�v��Ǳ���蛷 o��K5��U�D���ʥ(2𻝒M�٧@��@�T��F��\���V�[�k6]���_:�b�k/�������N>�~!@���<�����-_����3��g/����He���(z�Bb���T�����AbZ��
O�D���)t�ɰ�tS����$��gp[J��;5B9���>�6�>7,���s�7��y������Ӛ�q!�����.�����c�x��G�����O~ $��>�ѻq�Uk����}�v������/������g?�i��6ᩧ~����Q��u�u���'>�C��;��;u��}����ao�l�V�v���xR�|��f^BS(�HЏ����N��K�ό�^�r)z���^a��f(Ւo�BkNY�^-��xw&�RSB��Y?�@�\�LE����_�_��'�?	&�D�0���	7z�d%�Ölͪ9���*YEX�h�����͍&��nS
$��f������f���-832��D�@�M�)҆U��#�Ԍ|��Ί��Ҩ��	��lT������706:�T��S��4p����<�b��Ǵ3��P��4���l�r����ToA�DnFOU��dh��C�s\t��71'm���jT�*o6�Z��~ۮ+��n�B���jc�� }^�\����\���n���<e�j�zj1���0�f6�:d�Y���{%��6ꚨ����j��_��$�>4B0cH�:���
��\*�Z�L�ڠ�Q�e%�� 7�#�i�1�ӄ���N�Qw�}���#���vt���c@��l�_�1޺����PUm>G��@:�S��gG@AbZ��JѸ�C�Y9��;h��d�lk�K��-��SH���wR�>q��ᠦ}ɗ��x}:@q4J���H�?���8~�>�{@���FE�;��R�gT������S@�T*���7^����鳧P�R�� ����b��y���G�ߊ�[��� k�8��E�Tټ�ʇ)q�Z�عP��H�+�˕�*[�.Y0����e˘�Y��8146��h�p[n���Gq�� �l٢5mf|R:�c-_�W�[��h�dY8K��)�k�����6�]^�SYE�`�;�F �����*[��e Xb824,�B=��rf���S�羏��>v��Z;���g���o 靉��h����%��8���犺��X�\Fb^~���ꫮ��q��\D<����.�)6�	zc؝��C�L��!�p�Y���`%d&�n��|}ۡR6�����/~u��t�ھk��s���_r��ރG������H3y�I;T���bQ�i��rΦSc��s�U�B��Ϧu�'1}�V����**��XX�E�x�UTK��Y�r�Gw�ޣ�������������UR��d
�\�ݘ��U�c��/��/��M�:�$���x�&�ƧF:>'�9]�w���Ytwrz֮���^؉;�ׂ����'�u�7���{��'~�Y(O�<)Q���ݏ[�vO ���ѣg�����Ԩ���n��O��ûe��\���ǒ���v;�|F����p�v<
"�;h�\-��4x��:�4\��y����K�򗿢���H�H>����/c:�R7#C�V`�p۵X5z{�h�:��u�-�E��@og�f�ԸD�Z&Ww�Q���d��S���iLf+]?����	h�3o�2"8z�N*�.���]~���Ǳ���&cH�f���":=��-�����G�ա0O:G���0yF�`���SK����ު4gN��O�MD�N�6d)����^�[��i���B̔�R=��k����kV~2h�ӯu�Ȳ��G��M��U��K
�g����E�׀���j�����|���p�牛�8�,�>3W�$��ש��#���\y�djҏ�Ɗ_��	�H�D�UB}���b4x@�*k6�|,۝6	�5J�i8��f��%I��E��&Y��6o�O<�ҦD�~�:V*W"�%uc1���C�b�x��Yᚤ��f�(������a�y\`��)�S��J2z�Txmx_��[bu���5��4@tC�Û�n�BN��\�ժ4_J��
76�s���|N@e��=�I��#��J��IL��q����R��i(������x��ؽk*���Zv�_ԍ���ot��［�fz��&�b��Ы��6�d�8�9Y�|���y�*�{8�fȮ1�(!o�床��)%�z3f��Ǎ7oU6�>��{�nlX����P�J��M�ĸ:�V��G�����וןl~]W$�]���&&Mrw�%"m���{Y�@f���y���8t�0|��
5W�X�w�Ps1[跿��sӲ9�J��ֆ���Ũt��+����9�s<z{��ۊ�׆�6���	����X��н��D��@kSX{%����0��]���dr&���Hdr�t��������O���������X����;���Sg]�c#�������8�1o��L�sǘ�Ĥ��Ǎ�
�*��%�I;��HKm
}���L������V.�V�j�R,�k���ǐ��afj
7\���\�]{a��7q�}�`͆Ex��]b6�&���Ԍ�V+�q��;q�M��ӿv^�v �<��N|JL�����o<�06��E6��}H�j�lnEWW>�k����)l߾]h�b�>��c�?���h��~;F����j���܊�?���������SQm����ذb�c+�}���#౪���>�y�{ �V���&������ ����	�NM�$�MS�����ç?�Y
E��LiTvI>����黱{���E.hf�c���mA�ϩ$�F/�*�k
"B�]��:\f7J8ƍ�����9�L�b*U�t���g�0����ԣ�T:_��W�â+q���<{s��zLa](�����{��G2:��ێ��˘E��TȚ�S2�42"?�@��=�w��y��F�A��Z�k�����	�J|)�I+5,Lό�1�9�iWc{-��$�����e�y89*��b;m&Ւ�7oƳ��s3������'Y2����WK��b�϶1-5x%������h�X�Ru�h򲱡Khșw��[����	�8���{[:����: �`K������z'���������"�jjj��,$7NnL�,l��E���J#�Z�k^Q��p�(�R+����Y��?��T���36"���TS FH#"㸩Tmr�Б��ƒa�<+�l&�[�A��i��.�k<��{�M�'���I�r�kD�И�,	P�U���`׃���Vc���%���������_����;w��ɚJ�K�U~j\!�bkK�*ҡ1��ė>��<ro�|�l�n��ߎ�:��Ջ�M.�o/Î|-H�\���a�[��O�|J�3eV �H���
���SyL���Nf1�*b8^�=A ܬд�h�]�s���p��aٟۚ���܂�����Cڬd6�׫t깹iD��I�;�E�<8�:�������Vx��d������y�L�k*i��~>�|��y��?x@��Z �6Ηt8w���K�+�΁P0 �ӉޮN4C����R��ήn�wu+]��={p��1�'[n�Yz��'N���3�7�Ųm��5�	�Tv������˗*5� �/b`b�F�l�Z\{�ux�ٟLĦ������W�Q�V������V|:U f�	э���(p��0N��TU�3,�c����x��	���D��ቈc��=Y�@��!��8+����؁��^�[��"�46RF��D748�y�)�h�r۝w����4$t��-�CG��_��֭�~����~�ӧu�P\46��z*8�y�;eY����C9c�������>�K�:�Ōq?�{�=<�ҋ*�������݈ǘ48�Hs�Rb_�m���#x*���F�\�~5�����DG����J�������A�/]Mp�� ��ڈ1��"�m�m�B�O���9u���|�׿��#|�ŗ�(g�������\����)��TR<v4<h	�����cEgK#:Z�K�Ů���ٲ�$�cpb���
v>�<�6��șml��wzr�LL�a6�����R�~-���z��r��!�+��G5"���'�������+pxL3*�-�D�b���)q�5�    IDAT�6b�!���ܵ,m�N�z�+m�+y@�IuQ�F��'�'ݮ��K+�q�E��-��	~�g�hI#�jM��#J�NG'~.�N���:K�]
&
�^k���E��3O����\�dR`�iF]=.�4���(A���^��G ��v�&1�\A2a�1F�t�A��y�x25㚒Nu6�k���WJ'3.��&P��8N����D�66�3��f���A�mb+��M�-�jQ�(�39���%�k�[v�p�/fsb�)c[�_k������7��E�1(��X��Sdcm���D���a}�FcV�
f3�S�z�kQ�3��)�dh�e��Ən�~=3PTh\`��W~���{�Al۾CL�7��Q�`cuV�.8bT"FO��n|�k�}���?�W�m%ܰ~	6,�B؎����F��<|�l���3ʴYi�
)}fi���Sț^��+.�Hq�þ�l	��,&�iL%3:��em���i�B"[��tN_ �lQ��+W˾
��ڮ:��H3z:���v�n%��VK250U����Ip�g��_d��"1tV��-
Q���U0���0�6FjUF��{�T8�����P B�\B2���-�Jg{������r��!��X��d�rDZZ�&�x�����n��2�{� >�g�����I��H^�E�FY�ڇCA�%9&�^��?E�SnS�����/���T|�۾��w�S�/���Q��L�L�$�V�ھH�|6��5��oD*Qƙ��N ��!_� ��dZb/.H<8HPk����q�\8��-�
Q�|�*՜��lH��봡�9������ՌP��%:����G���#��a�� 5@ʿ�Ǎ�ނ����S����\Fsk'�o���p��i5zJ��T�tٴ7����(�
x}�v� ������a�r�JmԸ����*��x��v���+�.Q���{2���|ãS*�Cզ�1�q���ĭ�_��6����^@bj~'�;���ԃ*�c5���<��Z�*�	El��y\r���#sz��	���h�KK�2v�ރ������lT�}gw�B��g�'�d1��n��9F"Paϋ����JK�/�J����F/�w����97u�6I&8&3Y$S9��D��y1�v�g#l�^�;rJ/��ƅ�!1+�n<!.Z��C�qc��������3y]�ݲ=5>;%6�T� �1I�j����f���Z�&�IRs��4-�?W�y�ĔX�8ȴI���R8��*�m���ܨ?�l|�U<��&��ր7Yi>�߮t_9�^2H�"�΃hji X����Cx���^����,X�+D���;���DV;565��� ujf�䡐�/�=f����p2#��%+P��>�Z����-�ѡF ~�<���!;��xH.���&_�����s�[�T��,��90��8b���;�V�a���>?7A-��De��x���x�ϻ���fO���MC^fx�K:���l+N	8�SD�bs{Q��P����D:jj�&��bFƭ��g��60I���	�d��� � /�+J���苣�tM����d"��Bv@�I�3L���ѕkװ�����Í���㍽����/+ə��P��L�S)þ��0��nP���x�?�k�ũ#����ϡ�g�=7l���]hu���ʣ5 8�I=��+�w�{S�V>��5^�"�����b��s�rU�e���1��`2��T����٪��f�n������|�j9bCa�rm��f�J�ȺLL�(é"Nzz:��ݍ@�ڞ��sh�K{(mZm��v��'~�0�kM&��s���M!�:y��	1�|���7>�\G�I�WT%��r

���>�����kͺ�h�hGgO7N�8�>�6]�/�s/����[�o.[��W�DK�ScC(eS�U��r����Q�;Aa�xCM�46��x+׮+����|!�{�R@�R*������ Wq~n*�dk^5"-X\l� �_����"�N�W��7�wk�d����`��I�I�#�0��#�g4}B��j��>�RF-F2�Ta��t)�|`G&Ǿ��o��	��B�}&:cb�]|a�vy�bє���ꫀ �ش8�/�NI�Q���r(��Eǈ�2�ᥢ�4=���P��H%������Y���t}��V�7KQQ�wފE�mxw�d�c��+������>��Z���7���aKk�5!?��߿(\����*�A��Jx���G��+�`)Bf�g:�P!���(Qڛ	<*�U�@��D{c�~4{,��ф�z`��P�QlF(���阧�L���x�c�^�ʞf�iO�`�e��ఞ#.�-�����O�5ꙘC/��^���*Μ:����yʍ4Pɥq����ք�P�ʫE�\������3l�ZF`��g@	��J�W"���S��M�O�)Nڡ�!�I4�iKV�|�lR�4�,52S#��3�=�hLMGa�Z`ߊή���J�j�zܴ{��5���B@n<�l^�$�!��-V��').��1Ќ�V�5�r���Ճ�,(2J�My�hJe�������W>����?��Ktn���:�=�)�?���?\k�57|���H�����4\5+8O�|G�g�ŵ:���p�|pz���ȓ�ur=)������F{c3��5��e�Y\����Չ�x#��JR-�\5D���2����N�aAO'>��#¹�g��N���p;k4fD�n?F&&�Hg���a�GKt�T�Y��{�kW/ǹS'�;;3�bO�W�sCMX�a=��'����|��|��=�g_�&�B�G?�ld=b�9T�Q�T�V���Q���3c�x����-eq�M�`˪XSpg��憥S@�7@�\-��bE%��� ���
Ŭa���֒����h��1<���lc�ƒEL������UZ8����L��R���`߾}b��[��f$P�j�F���L^I�|�8%8<���T�6��F'6&��P�r�c��n7�{z$�'Òͤ188�Հ;���b/���	<���^7�*�N��i� +�XjI����ؠ�!?�#��o�x5�/Z�;�{�1����n��6�Z�?{����m�'�.]�˗�G[S�X����(�2�"!t����/V혷t����'Ξ���K
���q���=�ݿ|��˥���aTƫ����羙,Z�V�!N&Y9������(T��QM/z*�1�O��S5�
lbփ]TWj%��/f*����TKvYrP�&���cWؘD~���󹲀
��@���m���4�vE�ۥ��<Js�S�^`����	Dy!)�~�yg�C ��Fx}L�����SED�|9�|R;@�[ZƬ��r�{	](�tV.pN[_����нw�^�᝷^����""�x��O���Ac�>r��:s��s�? *嚓Èi�(���
t�����7��3�!����P���թ��̬6`6�~�3aR��JAm�a�a��Mt4���5��]͘�A13�\zNt+�8�`D*��X���%.Τ�ơS(�"蘷�=�5B;p�.�(��l��!Ҍ��݈�܀g�yF,ʲeK�я~/��<�FF����zm�}��[0��'����166��I��F���U�W ����v���qc>�Ն�~�t:�E���P�ذY�
\b�f�p�&�åE��6��9��U�F��LM�F1�d>�66ϖ5�H �;��d��-X4o>���q[073)�
���b�6��)�A&K&�Ip��>ikn���S"�� ��bzr���v#v�;Q�&��#�Nc2�B�Xd[���g�α���AwG+��:�bx\.Dg�����!�e	(�I� ��S(�]p��H'3F\(J�FAtoO�^�a�z�f''�>�P955���N��"�Ř;\ހ�#�b���I�]��[�ĝ�l���3�p�,��q�d�u���[�n��]o�o��{��;����u���(���f)a������:�~7�Gq��Y�}r���EګG��̅�>��f���\�IU��^)᷾�%��%�ӈ�ÈG�&1�*+?�Y[W7?���{N,����b����ܶ�p{}p�Q���Q|��t��Fo�K�t�뇣F+{�a�\�E�Z§n�7oX��=w5��&�5$�t���x~㕮��+���R�s(���!Gx�!�3E*6�+t� Cs	��XI0��!Y�!����W�htdJȨl��v	X	Y��?� ����I!i2����&ǵ���v���|�g�Z�+��q#�L��yj��ǣ����t(����sl�h���:uJ���8���.E�����g!/��^�X<	�%t�iD�d�2l�t-ڻ�mǏ�|w}�>,X���x/��������z��݁���J.�w�*�6���hk�7�_��j�~�����3���w�s��������˿2@������5��?��x��<�⪰:(�N�u1!EJ\�	T�`�6HZU��Eԁ
)e�'dV��@Β�&��M�"�,�T2�{\�+%�xQ�P�g���ӓڈT@X- ϗ�D�ik',V'r٢�d~� 3��X����W��].����5�.�~�j�\hjhD:KZ:����1kJk��E������VS�^  㩜m���1���}��{�q�U�PN�1p��\����p�wc��E�8�j59f�S���P0�/F�h2;�W��P4<yDg���羠,&P��✪��8{�
trs���S.��wv[��w���@ŋym!�����A%C�����4�����
�$	0K�g*85��s�(��z�MX�b#&&��ʫ;`q�̦��h�%��/	۷��W^yK�,�m�݆W_{��#��a�+�޾��������F�.cld��Г?7&�^����-V4�u�et��a�$��sb��������������e��� K���G	4x��%�r�c'��5��~�
����%��r�����Ϧ�X*�3/!�e3xQ�]�P�JY�fq���w��[��K�?��J�hcw�i\��ի{�ӧ����<��T0��P���D8���^���u�lR�������8ڨ��5��q��e�������������.G�6�_�u�V��M� @7����[�``dD,m�;w���l��&����i����Z����pǭ[
���!�ջ������126�\���n�N���([]�����}���{����£�B8��Ɓ�΁C([ �ۍ�kW�c�?}�U�����IX�!��W�X��RI�-%,���}��]
��ƖNkm�+�Z�2�"�^����	Tl.�L���X�����}(d�j!���T�/�<\� HWYSk�_�k;v��~����?{.�A��a���Ǹ��v�+���ɹ������%����Wʸ{�U�zI/Z�%De�=98l)�lyp�J ��?�$
%�$�f.K޸��U)����߬�W����&14�p,.1�D(Z��T�8K���S9*<���;q���lA[W��/^�j�*��r���0h���!�4�nTP��z9]|yp����l	Ľ^��S�&��HC�/����f4��^�K�Fd̘�B�5�:����ގ����e+S�Q�U�ߋ,<sT6l�
�P�?�/oߎ��~ ���]{���/�[.�n}��5�	�N��)��Ƶ��"ȴ�7��L�
螿��$�m�J�Y-����;W-g������_���<�����G�yG�lu�Z�͓>�ben��+��Y&�qA����l�^)+���|C%�9=if�es��`R��9�����8�A��GX�q^�R���c�?J$�q�R��Tؤ�L�*L�c�l�bʬ	v�QC���I���*�0(�$��7Z��� ���Q�i�r�"����<7�"Jz��:�jI��r���z�����B�j>k]MLwt�����{��vভ[p��͆�q�8Ѻ3��J�S�XUϵ�5Vܶ4?�#�+�I����o���i������@:���/�+�3�(ɭa�Ҋ�h�3@ŏ�F:6�7�Ĵ8,xl%�f�@�,v��9�2%��v��s8;é�iX�-X����x��dϽ�MVFR�v��
��ɇ?%��믿�~&���.?rN��U���W���_��ϟA>���IƦ�����pC�@���EN\��v�̛������L���Ǻի�$�,s�4'PǮ�nQ�Ǐ�F��g�]Ru�
����Z��52���_�	֭��xfrR��ɑݘ���L<�l����"��j��IO�j����mX�h!~��_A�����Ә�Nk4�M��N,�@{[�Nw�>�.����`8�W����v47�;o��ZV� �a��b�*+������^;}'�]B4��?F��UYy��ʨ�S���X�x�/]�������'�-��׬���$v���BMm�reh͠ �Þb�z�.�=��\K�c�"����-4DhAu�����?w�m��%"�s�Q�gPʤR�ؽ茄0p��
NO���ɹ�JL:]�~^��2�x�im.8|!X�Խ8039١|V��=wm���^���j ��0pyH�Z��N���s���
�W3ǎ9�B!��j7�p�ޱB:���-4ٚ��)�sY־y�Ѿs�.�����;�9|���1�ͭ��z�ˋ�1*��+���o�XjX������G���el�y�Ky|�p��U;�@q-a�����,ܶ���,���t2卅]�Ӽ*dŨ�"�R�+�"Y�b:S��l�s		jg3e̤�PS�n<�0FƧ�`�2LNGq��Y�}�=��3����%t�w`��:��6=���#��)Ҁ��^9*gf�Ō(ɖn:U,0ߋ��M��ԛ�\�$$�H�Q%�佐~���ê8܊��������z�Jtuv�&'��T��{M&m������+�^l��&�}�|������k�}�[x���06>!����+�,��aE1��Fjɢy8b���k������"0:9�h2����?�ޙ|>�g����X��/��BF?Ԩ|���ߜJ;I���\�"*s���/$��@�3F���d�Rq$_��bэ�[ ym8�!�l�������2j����d`�ZP�G����,��v+��,b�9T+ti8E�����D4)�.���.	��lRN#�97�NP�� n0��!�%V�3�]
�q^L����)��c����9���S���V��΍� ���F�a?海�^*hNf�h�����ǂ������h���ȑ����tL�٦iG�`����H�@��u"���"���^�����9�9y��N�Tȓ׆�q��ʱ�6G:�d��f��jy�V��Bg��,�.��\hx�c�@"�CR��T�R3�<�D�VĲU��4
_S��_��.���8�]QWI��v@z{�����ʫ8v�����C-ǎHL�㨔r��g��e�19:��jfj��/��o�F�C����R�?�:	���'��Ӄ�~���$���r+�/����Z�9��R�����S׆¶�����A�;^�*Y�*0��T������r3B>/�n�jߙ��I���e�={�"�+Xlxc�;�i������d�r�VW��W.]��kVK�R����r��`zj�<�Ex|zZ��sP�ވ��.+��8�h�k�?�ɱ!� ��,&Ƈ�@��X�T
=��Me����pB�v��fT*.��K�R.��M�j�B\:s�؜��eSTmO�O��n���.�&b蚷H�G����ks���7\}5bS������a�O�d��#��X�j-�^���q8�a�)֯�t`*1�UV��荄	x�R$����$��8.��x�����}�"U�����elj�h�c�H`��Mغ�z_:�s��'�2�������8p�$�\�l2���.�9�u8ŘT�Р����\#�.�1���0Aj��[0��sR�{��+@��?��~�������iT
�:E�@�8���$��[����m\����|S�C���G4���o�`ӺeS)�V    IDAT�f�R�ch�T�쫠ўG�VD)5���<�,��7S��8�t{�&�p���*�0�bx&��lc�$���Ȗ�;�Ξ��Џ&��n�t-FF�q��il���I{��EcC�BM�'�1���G&�՚E#E��r�٭X�`��6�3g����-�*�ي�z�K#�Ѷ�MO�x�R	�������кH;:�認N?������l�/���	��v� ��i��8#�+��BAlذ�ݝr5����~�k�ۢ.�����K/��X4�}��ܾ�.�h�n�S� P*搜���%���#Ob:�D�\#�8��x�D!���?��_�r��l������D��p*�f�vX�v��H�95��UA!T�
r���5����r��`M=�I��j�	�tK��"m��*եb��B��x:�(�?.�N�2�d.�+W.���N�>�|��#����ju�4���a�VP(���:l^	|��ѓΟ����"CcRB���7��(�N���0R��Ҵp��¹b�X���_��k)"� �u���m��� ȋd&��k��p�z��M�6��M�)E3_FDK�͑�0b1�dɨx<�ͦ1<<�s��	��^�|��9�gΜF*�I!�M��$��{ɗ��	%"�q�8��T8fGgď�F'�F�s$�1��6��ti�*���偼Ճh��b���)�t�C��U8t�"/Y�ޅQu��p�Ҟu�F��ؑ�8}�(f�������&�F���Ӌ3�OIP����b��%H�g��]�x^''ef�H��hni�c��а6�;���<���b�8���n��e�m�-�$��,��0;7�?��u�awbx|M-ݢ�9Gw{=:��S˥�P5G���f�K%���M���сTQ��pit'/\B2W0��|��-|�������.@۵Aw��"֯]'v��R��3�.�={qq`U:���u�t�cv6�¦5��ا>�K������Hģ��l\�����/&`�����n��*U�\?t��ō����되����0.�׉��A�ˣB=n�t5:v
��<BͭZ/�t�+�z�N,_�7m�c8s�����O�	�DZ[���ى��)��@c{����G�t��{�z�|^��g�%�ĩ#�H� ,��d�&j�����Ri�� Ó�pllB<��M@��ۍ�7�#�ߌSG��¹Ә��R	kc����tt����{�ݏS�/�Y�M�ʞ�p��0b��n��69�N?"a*m����@���0�d:�V�RŊ�}���a<��Oasy���"�Rw_R3Ù��cet����!ƃǼ_�����3g��?��Ύa��زy�\h;�a��A��G1�����d^	����e�XߡQ�M�\	���&Ee�L����#�/����k����czvVL��<������Qp�w܎}{�bjr���lF�.�-�W.���)���(&&�toi �D���T��-����q�@�vx�K��bl���E9���q������(��K&��e�-�Ғ�]��a�W�DF�!�iپ�t�b�D"W�롅��P�D��S�eտ��b���� ^y�5$���c�LF��ED��j}�3�?o�^/�hDHзd�R\u�:��w��D|��}ﯞ�Xj����3*g���O��㉌��t���@�T�����1>�y�/��x"%5F:��j\�y*4aJ���i�J�H���b��~FwN�|�2��D�堛�cn��b�����|���q��AQfU��+Y�/�P�z�K�����t\��I5��'��
�ZĿ�g��婞#��	H�+��fEl��LXT(��\�b�4�����p[�j!�;G@3O�^�f&`sT���a�Zl�z���8>���w<��Q��n�&��ؕ����m������u£�� ���W�ý�=��t���i�h�9��ō0��\h����Rf�[s�d�0֙�VCs2A���˃�XJ��^D3d�\G{�B��\�'�{Q�@_�V6�����Qz'si��$�.����n��&�?R0���=���4��vlX�
�T�x�TR�;���>�f�#�T��!�ܤ��Ҷm��f�� {�q�:<��#
��sW�她"�"�x�~�}�8z��?��l2�)��#>*�-�����iO?&�h|vӓ��.)�!�\����ieoHpK᜝!pV���H��G_w��<rٔF����D�L����G�����ޅ&v����ƻ�v�W�DQ��sǫ�c�2*
�r��/WKdp��9-��66��bq�=����cú��i�U�P�:73���	�}�Pn���&LM����s��	_�A��w2$9ZC�9�wt���X��S���K9àV�X�h!���䳗10:��P�M�b���F���nŖM�v�B�_���Oh�Lq(�G���2Gf]Хs��%$rY4�t��Y<���~ê5x��{������"���E���X:�ff8q�ľv��-�SM �?�y�	\w�f,\0ΜV&��'G����V�A� >*�~��x��	��'��Bق�vø�Z�t��h;��o�K��47���I���#crdO���uؐK��v#vc��~���h��������
{��;����\���+T�b�v��Y<��L"�\�!}�x,��h
�lpx��5����Ĵ��J�J>���48�7�ܥw��_�"N�<�ݻwc~_��o������ϞS���S ���1�w+���m'�S�Y����vEק�it�uJ�±c���=�d;.I'Ąk���{N��b|6*1x6O�·T2�kK�/�[K��z�){��#���DB��JsQ��?��X�l9�}�}��O��Z��J��n���Ɔ���.��LZ��,B����e���1�Y��r�ء3�\�[/�����W�HL�ԮoOe��q��*��7srE��z��EX(���v�5Ba#Qi�T.��%Ѻ�ԩx橤���;h�%Be�����0k�F{�ͦ�=)s2*dU��.�46q�֛���ށ����0;���L�-z^r)��m��h�R�#ɩ��D|t(��嬉��Q,V4\��5-��&9
��L�G�����Qe'
`c�F� ��x�E���h�p3͕n'r��Z�7��z�,��L~Y�t���ϦL�9��\rWMOGq��	�����).^�]w�%������X�tF�B� ��ƴ	���{JwSg{������٤��F�熥�G�焗�;��b2���c�5[pqtJ���w�}��ֻ o8 kŭ�p�t=�4�tY3r�h���b��E��g !Zxw�^���H�t��X�`����I1d�u���ǅ��q��	�Y�7ߺ��VQ�?����R	ѽd�l�w�v��%�E)�Cjhd��i6�ȉ3���D�Fy$f�[��ٕXL{�c�<,�u���*>�F�jt����g|zF�_�\6Vn������#�A2�sJ��l�"�w5K�516�l��?��2kSsQ��O����.wS�4��!�K�i
�;�Ңz��LOM�^@��E�2��2yL������Í(���`AF.�s��kt��(N�8����e����VE�7�"�x��`c��7d�d�/09>�'�Ba�r�uʢ���ts��Z�x����/�1�@�Z�\��9�N������^V-],����X�v�>�9�8Ć�9�X�8]hhm�)?��c�[8}���Epæp;m�|�:;ۯ$�R��ōU�C����&��.�>����Q���^�
z���҈��O���c�ho�5�7Wm�Œ���`󖛱}�^<�/OI����'�¤T��<hTi!f�i�P1MԦ8��O~�TO��?�0�
5wĢS����Z@�ǆ����!tGB��@��	�$�Nf��&�造6S(a.����O0��!O�ӃB�,kx��P���O|�/^��/:�֬Z�W^�v%�> �VEg�漖��z�N�&�}K��ۭ�Ⱦ�}���bA"C*�կgMuYe
h�V���ϟ�ѣG5v�=c #o��	���K�`�r�=wAf�?,֐מ��Tu���L!��H>�*SSҵ1��Nˏ�X�jΞ=�'��rY4��3�z�jE�U�ǫ5��
��jlL�-#���-��\�jY��c犙ط^��_��b��:�_��/D�2X�6|�g{�=��>N���S�j�-M�{U�Z�G.LdV�3�L�>���ev�,{�
��QQ��P���,���fy��؆����E��T�~ .X-n�n-�#~�<--A$�i)�mv?N�������جN�,�'��ثr��t,QY`��`A)���܆�F��ܰD�BTn~��B�422�b�xr�5�gb*æ�aV�y�n�57��ZZ"H����؆.�o���n0�$�J��F�1��L��	�2X���~�m�x�MLLM�����1q�#��X�v-�ɤĥ#��q�BoMn�p�FbF_.��x*���%=88���)�#!,�7_½�ܔ�$�D穅"��~��ܽw���y�y�|�N��9�4IM�I4 @�BIXђ,$Yad�z���ge{���lYX�
����&��MӁ�9WW�:U��I���~���?���;�����S�s�����y���W\��V\�׬�o{F�_zMO]��i���s��X_�]���4!��Ď��F��?�IM�<YG��om��ݻ<bؽk��.��K�_���&�K4
��;�����`��z��>���)޸>lntQ���M������w�!�SI�{���NSsk��N���gҾt�&w�|���46:��ŊK/�uyc�g���;0�C��j������}�A|%��	�uup�^�}c�6o��krҬ�:u�I���G�i�i�<��h�,Yb_�8\
�b0�|�����K�5�2T�����7^?�}��Z��T�s�yF��&M���VOϐZ[�������~i���S�lX�"��#�wS�Os�!��/�H����|�1<+t���#��ǟЛo�n�y�g��sϱ:wXPQ�	�����^�3�>�^*H[1W� ��Ss�E�>���{�ib86�3�,�I�f�g�;�b�h��{s�5W�s�4��N�3ǅ��H�{�`o�^~~�^y�%%je�<{��X�
S�/�����-�|@�fϱǉ��vi����q�ݹC����:|���:���O[��(t�f�>�[-��b]v���b[d����m���a�7u�l����aoF�e@Q��A���'��1}�#������޷�E���&t�!US�4��ZI-*����.͜ڭֶF�1�ō���Z)�LihxL\�	Y=u�D��K	�&(W����=�Ɍ�n��ھc�֮����׿[GҪ'��g�
��s���Suh�70���י�����{�N��R����t������(-��h~X=Gٯi���:|���9�4A�d��(�oρ��->y��:��/پc�������Q`4�E�(�%��{R����b��# 9|M����m���f2��.ߧ>y��0WJn�ә���|��Y�tA� !4���.a��ŚwҬ��-뷕Ǉ��؏����e
�=��_�'�h���4Z�=��2x1`�Mq����,ˌC�߹)�}�p	L�'��9QAA��(H��j�Z T#�d�����w�d �֪�J��h�E�.Pg{�Z�5s�dH�ڵk��ҁC�z��:tt@M�6�fc^���h�K&��D�!d�~1��46�|h�^�h�qE��@k��0�&pu ����w)o�.�2x&P�� ��;�oFGN'Ϟ��3�*�����!�C�l�2͙3Gs��Uc*(�J!�q�ˑ#������7�Ү��u��a#A�IN=�tM�>SO<��2F�#ǎi׮]�54x�_���Ŗ��gݰ�)R)T8��B<�c�Ūe��3I}����3���@�vmw�fo�]v���`��Xv�6�ܣW׼��[���s/Դ9�t��i���;ۖC1�]�x��`��d�a`ӦM3�2��C{��������_W�A�E�F��y|�sh6p+�_z��&���Ԓf~�E�*o�]gG��f�sX�Q��h�#k\/F[KN=C3�����Xwp�pP�dJ�ׯ�,������ԩ���*�Z��לI|z:�ɪ:�9IM-�&��*�W&|:�O������G�<��x��GT
��xA��.Q�R����<����՞=��s�V4� �T��)ػڻB�@1ȓO>e���?��o�g=�
ep���DU�v�Ў��=�"|�g398t��L�x�8(x�]S�j�+y���=���w�N�	��M��Y���0���)��̛�vB�
E��"�qs��{�u�F���SI{�̞>�6��cy��G444���e���
�����@�JA�8�?������5��ˈ))᱙��HF�<��F��7M�����+��%�F[K�_���(�#G��a_��"W��!עM[������Q�kf��xp��x��L%eC�P!/��~e�\4^�.��Ͻ�j%6`"�Ƹ�ܔ����]*Q�<;dMe400h����S2ۤ�y&g�*@���g%Sd-�� ����Oӳ�=�����ӌ��u���T��D����i��@��[�M����C���O������a��i���SO7�ƻ�'e�޶�o��op�Wccyt�p��56��vbxh�^B��St�+�kj�����ٍ���%���Z�D'%֌B�6����gæ�Z�h�Qƽ{�G���HQ�b�g���LC=�^���;�����5ʏ��Z�ڎΎ����o��c�(���RyG�]�Z��x�k���X�
�z��1#Z>����Rx�́�^=��X�X)�}@�������J����(T�s.����@-��5;i��g��Z�ʦ��:e�V���G���F���ht���k���6����� ��E��������
h
E\�&;���S �>�A�n�!;�]vd�`)����2�Ȕ�QI�}�.�����(��e�y;���:)��tj��LSkG��r������$�}�NC�G���70|P&��4�'�n�G����t��A��������S^)@i��~0!����3�`�|�[�n6��y:.��=7h�E�����T���R�d!P�d��1I3瞬�Ѣ�5���Y�.�ɋ��>:�T�#̭0+��"��Ժ
�C��)�z#�L�qK~�� v£�2���P8т�[՘k���HP��J%�.ZY����K%l6��5 ?��!k�Η59���>�dF�A̵c�p<tȆq���V:��c���ۼ�@�e�#'��ґ�r�`���ؐnP6רÇ�<%56Q�FkB�S��ʐ$��/U���:E�L���AmA�:
A���yD��fΞ���	�N�H�Ө:�t�
B�oߞ���R�y-�C�����1M�:ͯN	��r]�¯Tm�H�O�9w�,���F�Lf422
�uk[{�Ǚ($$?���V(�h����Cpt�E�j�V�JFv�paGw�kk�s�}���⠀��:�GĈ2�csm&��%�\��!$�SS�F�������샔�G�97�@���5c���x�P��TO�Z:�:[���;��k=��� ��=�Q�z����fLn�g?�	u5���C�s!�2�T��L���-9�<U6���e��#n )����b��(_��}�:x��f�:I�\�)�C�B�θ�pԙQ<����]{v�gV�ءC�=g��bM���*ˍ��_h��]�.i�^�G]�"�y�,X��7w�q�8dU����������ر˨���;L�E���C���ȀU��vY��E�I�&��	���p���\�d�E
�4�<o�����}����)��"�?�/�m;wi�}ޯg�9��1ϋQ�$����'p	i^x6A���;�~�� ��T��<���w��yw�������G��J��ޱB��������k/�s�x[�2�
�� 9�8����@#0�ˁ�¡M2�y    IDAT�Cι#+�r�(���m~�`�y�,/� 
Y?)np4��)��7(�Д)�tǇ>���׿zHcT��&�S�FUjHx'̴�ZvX��jk�M:?�-�J[s��v����#ajtJlV&	��t~�����
�C�C�U9׉y.\�P�a1ݒ�)U��;MR�t�:�E*�Y)uϡT�p�d�'�E�qw�i��xMT�==ǃ�"���5�y'��d��.8?�h6m�aE�
�&F���y'�ޅ-/�j��n�7o�fT	Y�����ZU����85��Q�ɱ��=x؜,V�D-9S�|�!+Ktl�(^ $f�I���������5u����PP� Z����T�$6��v�l�NGD��]sǃs-�����{���C7
�c�clio��u��?(�}�I��/Fl������3�z#��10��>A���6�$r�1������ ͓156"������q�Q�R�PT��ɺ����C�|,Z�u���Hq���{ �GM�</^GGW�ɜ9�m�19Wp|��{��a#��.�˃�ل_�>��?��{t������^+��l��wO�tY'�s(�(��r,��9����9���̿���"
9r��&{�P�d��,��Za��w�O�	�xM��3��Xq�X]j�B#B�&ww�+���)�6Ed�z�����6b��[��t�;�_���
(܋/��}��3��}y��uA�[N)�m6j�>i����(����+�\�xL��L5A3 8e�����x�B##�{��1*��!�=��>�g2�:ԱbuS��I#p���4>:b®��h��A�_�Hf��Ƌe��!�70�*�3�P2m 6@ɿD��:��B���ဪD႟�̧�~Q���� qva��Mb��io���{�	MꞢ[�s����o��f�G�xa��n�w��4�v�1�F��4Ҩ�)[^Pb�GFkԙ��51;ϸ�9����kR!�|p���TCM͍~6ͅ,�h����m~bt�[�A���1�F\(���K֐��溂X���EBY�d�wޜ��|���~�=+��_�P�Q����K��w<��|5�2�d=f��h	&꟔7(���WJ���2DuZ,�%W�t,l[[�δ(��#YB�d�Rۊ2��' #E�Ǭh�D�cs�	%�WB`w���r�� kּ����R5a8Ń��42��U:�e"H<!���m�F��܀Y�k����=�
����8����\���	7Yt�rA��0�����R.�!^V�4��H��;Zt��3�`J�ơ}���a��K��/�C���w�eqͥ�;1��s0в�:p\ }��i4�6a
>��{Of���B���t��]��y�U�w����7�	TS:c�#�K=���j<e��޾!�HXO�-�Xg�u�~��Sڼy��::�G�ω+����5��%:�K�	#?v��2`�KY;��ݪ������;�"�q�]D�\z�ud��8*�P<���g���#���)�)��'��9�1v����N!�/��h
c�2u��9�{|	?�~i�N�A��O���%�[sg϶#/�t)�	�PmV��,�1���N�����mX縊p�T�o$oc���N{�Ua/�D�(OcS���
y#J7n��oo���c���'�Ġ��]"/��4AE�GX�^k�����d������⽏cNa5:j����1���T����E[xulI��G]�$��J9T�󱗇'R׃��lWX�c���H�S<�'�
^C��M�R�m
Db/܀�8�BA�C�^(q{��t�>��?V*	�j�Q.�4���{~��_�[�����Z��j��^tх����[uww�+_��_���E�ص_J�mD�gZ]����絃fr֏+n4��;b4�(�����J�!%��p>Sͪ6�Ō�cRW�ѼfL��_����ScK�k��(
���
��Zz��vI~��W��+UA�*FYy�B�$��!C�����&��a�Y�p�����w�g=p��u��aM�>���xaTyH�<͝5S3���h�m�3w�>t�ͫ��}LPY�r�|[��䞻�e���J��"���L+�z�Dd��SMF�L�s���P���^�*�0
�����q��j(��~��Q�0rwF[�IC�_oq��ȣ	)?6<�(Ȝ�ͺu{���榱r1^�t����ۮ��sg���;�yG��Z��_�}�?-}"��h��_'[�o���X����4؜�>�N;ӧ�݅���9)�����Ma?��ʑ
�$�P,4�Ć�����#��2��b��֒2I� ���d��7�B??^R�8x0�U��G���B�!dڔ-5�����c��A����>��7w�A�	�6#f�l n�,�8��]5k��2H�y0�ihԘ⥼���{4��YK���U���?��M��0_@�Ã�[*��U��OySB�J�,rK�Et�~n����B�h��eB�$�A�D��u Z�d�y��y�`o�k�.Ɲ�a�p����� Ƕ��QC������X�w�����."�G)
�:*G�ņf�r�v����Q �E&�8���?�֐	V<l4)<�(A�kD�[ևE��z�·�Q����Xg@��QK?��8�ɡ��=�,�(�
߀J ���}Z�I�����+x� /��⋵��K�B�����jp��
�yX�E:�t"� DPJ7�z+�gŨ����M��]���8��꼥��!���fLt��e2�=��cEQ:�d%��3����k��in�ܝ��J��`���$(H��'ൕ�6J�ڌ�S��s�屐��H�Ц k���|�$däf������\�A]ث�U@~�H(?�ތ��r�p!���̏�Lʸ	��!�*M#Uj��bO�˂�J���F=�ۇ�i�e�����`=�_���җ?��;��ۿ�{�?tPW\q������7t��t��7i�������Wz{��3�ǁ;W��Ɍ;1D����]�h� pIsyX��+�Y��raT��Rt�ɱ�0��	i���?�Q]w��ڵ{����-<Ņ����}=��a�t��;�k�ɧ�X�'?�W���s�'{k�{������� ��)��M9�����1�w\���L�_~����}Fo�~NS��V�)�*d� !=y"�#�j:�̳t�mvt��2homV�q���h͚WUƿ���2�DVq����(H���µ��僓�NZQ�U���Cx�G�x�1:���xd�@��Hys@i���D�
χG���[��W"R~���f�r�yuw6�86��ژZ������ϽņO��w�P��_k}pՋ�ۑ��'F+��zasᰧ�`#p.�b1r��y'}6.,i�Vќ���ɢ�ÿ����&�
��J�$�f]��o�3�� �%��#��c�C7K�UW��)�29Cm�@,��������c�P���X�>T���joi���7�ё1�0/��-U���9%��S�,H��!�r��.r<��1zJה�
�2n~��@�&Ɔ���;�9`�	������&\g�Sxp���m�6Q��pQ��>�6J�Ru{t����EK2��L���@&C�G��Lx�>c�4m۶��1�;j�K�j�z�БX�7�7R�ܥ*"�D��ˇt�a�>�3�V,`���,� -	���2h6�1���"����ޘx/�f�F�Bk���M��%�r��aבN��R<* �ē��F.Za{��F�Q2�O�uEj�<#PC#��TH��͹����0���Pݝ��ɏ�ޞc.�}�jA&A�B��gS�0 ��,+6n�w�Ee�A�+�U٦f_�"FJ)���m2�9x�,FW�}�-Z�j�#�1��<i�I�<�����E��3ZE��A���
q���_R���1�kMghkPN�N�N��i���'BSqUpĦ�wC�ה��-�D(�t��c��bd����da��~h(�2j���&K�����P	�-�R����z�O1�ٺ:��-t������w���zs�^#]x���/�w��q�FG
�b��J�Z�n�������W���7߬����pH�'Q�uOҟ�ٟk��*�"�3����z�	�g.T(X�� ��v���aM���\������T�G�:F�3'M������
�[���谺�N��]�ݻ��'�02u�����[�����˯h�[o���cF�!��|q��>Q�2F	#�0:�7$������zeϫ�3��x@����8m|k�^_�jM����,9����y�]w���E#!m�-'\���ٻ��������htSl��'�'��K�͘��^�>5�M���AfCSI����^�>NAl�:�1�EAE�q���p�ؿ7��WE�(s�<�(�6�������C RV�P٦���\�ٳ�8��}���7͟O��;��*�k��W�<����ʗ�-]��Q_����LR�sP.a��A<<� ���p�uq�""�y^ged�$8�|�#�3Dޓ�
� ������Ax���ِm�C��55g-��!����F�z�|*W6n4��6�`[�>lT,*ȴ�86�̲Ӷ��
B��
:$�Bـ���钑��$����&�y�]v��X{���A4��je^�Ԕ��<�Wߑ��+���/�7���(�)Ň�3�1��=�`�ȃJ�́���idǃS��g�Q����MO ��xv(:�X@A�-9 Ъ)R���f#8t�N�&��ݟõ|m�mܼ�sl`�r�\�@���5�1
�>1� �Ũ�`d��&�,�l�L�#��6 :;PFf����W���65�b (�L�K����Z7*����뉒�%�!B#}d=����h��q�_)+rL�P6|��؀�{j��jeK�I��)�I����"%��8:���a,�$�!�w&��/+a���4��c{�d%�mC,KiR�%��!@���:���;�������˯��}��9� �u~��k��=F� �^}�5ڲ}�ּ��כ���Gec>@���A�Z�ڼ��b��b%?Q�<yj�G"v)�w�!9��:�:<-Fl f��GW9Ȝ�l$��CPQ�KU��҉��"�<��[4�z|��z������0���$Njx46��z7e�S3�{L�^t����;�O��=��q�+.�H_��W�Ѓ�8���WZ�=�)z��_�r�7����׿����]������a�v)�"��)�5m�l��`�o�6ۀ2��RF�0����W4:p̦a�]�ùȤU��}�5Ͼ>��]����/#{w}�.��P=664�b_]v���>��g�s>M�
�����͸8���7rx���`,�ƈ�D}�L�мZuV)9����O���g�`ݛoh������a�&B4��5'�_�ZZ�����'��~�I��cV �솂!��"�>k#F��TT��|�E��&��D�g���,OS����c�}z����-
hI��'µ���Rts�x�a�3w�2�&��7�E�8���ѩ�]�����o���+6,�4)J}�
�w�P9\�5��uk_A�TI������XM۶�ӆ�;�/&�ɶi8�ܗ<�`��<�J���
�].�GR�Y�叐��$���lc�p8�UtvM�q�+-Xp�n���ڽk�V�z�J"�u�b�{9o�:���t���C���"!���^��8a������z��ijT{k�N�������;��^��a��E�K��a#sWb���ϸM�X"%j�/�1�V_%c5�jJV+*��Vbf�d���t\�b�h�/�@�u��;��\>Z�Rm]�@d�ɬ5�	�{p�u�@«���[3|����	@�4RK�+�1L�H	�=
�fwp.@WlR�M� ��W�΍ၥp%O	;n���P	�I(�N�%挄�����x8,(T��Q��g��d���G6[L�8`,)���*l����ǠN�4�ϥT���k�P�_B<f+�F5ؘ��A�%~sZښC�E#[r��wfu�������~���W��q�9����,M�m&ؘ�R���{T�W�V:Aڬ�ԃ���{O�82^�p��\{�[;�i��D�E�%����{�?2���n}��l��3���y�\�˯\�����Ҫ��GZ�n��4W_��W���/��|��$D:{
G+�nLXN��� �4��8ɼ��䰡1�T�2���@�9�"#\;*�)���{��!KKG�!��Tq�"%j���B��pH�B�Bp'� *pT~_�x܄#9#F���DΌ�M��#*_����vmް�c�K.�D'�9I�7�ٳ�j�ʕ��7�Q�s�V\z��n}�(�׾�5_����6�t�M�򗾢=��?_r*3��Y�=�rM�|�_�G�!������:�;2|T%�QnR���fҪƫ� �����������_��o�o���Ȝ�TբE����?�%��C&GF>�_?���\�^cH�3Y��Y�4���q��є0��bl*�7��~?>�d6k-�{��Eꒋ.�}��ؘ�z�e�F�9����$��U�6��6��F}��KGt��{p�8=�8Ƥ$G#�(�w�YqFc��"EK�F����Q�g�PU���z��
�$MHNQ�>��S����3�`+\+����W�Q���1�#��M'��쀀|T��u瞹�7��|͊3��w��)Tzj����>�����w���������Lױ��~a����x�&�a�����4�p��28M�nP����N��E)nt�:�p������OK6ݭ�읟��G����&�N��*�rH�h�����詘{����SG�G5n�F�2O� ��H��A�3���0�y����3���^?C�#��^������Q�F:�E4��~-�u7�T��y�l��R�U���DI	��MT��L��9U�R�p�qM�+�M$�l~�Ȱ"�I���l�0���3�J��q1Y��/'���h���P����h�^	����ado04c��; ~F�C�-'3� � �+�ˌ�`�X���3�zHR��gI��+<��/ah���Z���C��B�*��|��`�ļ�%����ߗ��Bȣ% �d(2������9�&ѷ7%���'i��I>�ٹcGNL�ˆ&�M�F����=�[�X,O�s�����{�Q[[��-Z[�1_t�YJ�FU��8ү��~���i`�H�T��88/�V��MȌl����5���=B(�SJ5w(�mS��K�#%��50:��[wy4t�G?a���5k��;�`�����Vi|����{��������|Uo�K�|׿�X��)���f���l04���-M1��	�
|��vH��<�𘌈��Li
(P|b���q 6�C�% �� �h�!�~��OD%Z.�-�Fd�
x�0n�8L)T<2e}%���g�X	_����V�S�5e�:�sDO����q=�����#�խ�ުϿ@_�������O�t�|�?p؅��[���;?��N=]��|]�7mQ���2fY?�1k�u;:<�*�R�"#�h8ĊH�SqQ��4
����2	3BT�'�l�4�[��O�B�ޏ�V��̛r@�{|�s�׺��i��m��Y2u�t}�����w�%��5���@~@���D�@x��@�g�g��a�p�_�d\,<e��͝����G�4��k.�`����	���h�#"	�ٳG7������Y�~���S�������D�����5QDLD��3G� In`�'�	��$\T���n�$���o�7�bѐ�n�>c�
�:�m�F ��Y�5BN�����x������b�������-�_|޿^�r���.���S�yr__���u�~�����t��ot�7��KpEl�/mҮ=�/�m�a��#�d̤O敌Q`�{�a��r��M)K�_%6���sfZ/�C��{T�6��������st�XQ6��x-�}�鵗י�9k��u�jojQ_/�r\k��-d    IDAT^y��M--:묳4eZ0I
�$�7�Ё����O��w����,s~
HFa�h��]̪g�ӱ����R)k��Yz׻�V{'	�); ���Z�AXX���γ��T:�����T�TV?��6��K�xZ���E�jF��T�J�J�(Zb3U��94�d1� �� /��<ٰCRu(T�����]B�9D����:a`�b%Rd��S�x�Q(��9��Z6Qa|vx �p����:L�" 7��ƥ��|�1��j]`D���U��7lc��8*�x#O��{�Ey&�GT��Lʍ�|m�G\BPp��if�v�	��{E�#�����ᐬ��l$��80n"Ǥ�2eR���b��.Z�q&�&2K��־���͛�/�ѱ5��j�͖P������F]w�5jH%��~�L:�S����^�%�h��~5��U���0ԯ�h�ҕQu6&�֐p���o���'�R���6����4Z��7_ҸҚH4(�2E��i:>R��DB��j��ú`��:x��v<��~�s:60�����g��W��ew�/����-;K/���~������0��ۣ���qTX����a��~:�$��&|�T"����=�U6s[�G#eȸ�F�L�����Asg������q�R)�gcGg���{L&�֌�"ycPg+J�b^�|.� k9t��$�/���c���K�������_ߧW^z^�㏴|�yz��t����y眫��t��������h���?|��1G��X�>�'�թKOӷ��=��Ǖll�8�Y{��P H%�l4*<KaTA��B�����U#���"�7�k�P�4��m���������~��r@��=�,_���}���뱇��g�U_o�	��}�=��i=�j�FF�B�@ܣL��K�9�&�g7"��\��J�SU�!N��j(�� (�����1sg�ҔI�hk���Z!�&���K����Eٵ}�	�A�g�b1x8E{"/�6�ϖmJ�T�������R˒pTbI7�樀NG������ۊĲm@h�Al �S�P�x/����V�G��B�^0�ZD{\�6�$+~���lV)���XL֊;Λ����}�C7^���;Q��#�����_���+���3���ы�_g�.]�R�ZZ�?���W"�
����|��EM��ΛM{l���R�B�b�N�K���3tޙ3�xy��#vқ:-�W^٨��^���Y�gw��xE���+ھm�x�WZ��|]}�e�����:���i�v�����0��v��g��IS���-2���A���s��=�F8�0"���'���?��U�Y眫�чO��ʫ�����N����w��_֢E���;?��N:����c��������mئ��	�0R��~���Ы2�)+++�H��"���U����x�l�X͆Ku�����]�=r֦`vI�h�l���CߐbP���s�+�	�Ҡ��b���L�a���>��t�b "c��������8�޳ZU~tD��@�5na2sو��J���͆�2C1f�!BL�����,?���	� �10,˞cG0��T�����p}f�&<��� �Eh�*�7�;��d��5�ܘ�Gks��=�l-;�T�]��vn��8��l(�y�N�t��z����Z��[n��/��~�+_k��Q
:��>�K�6g���}F���=�_��xQ{�(VR&VQkFjIV�KVԔ�(+�ξZ�qΧ��Y�	�!�?�ݴ����+i��T�hU�jZ�T��y��ۧk���Ͻ����ڵw�֬ߤ�~�NųY=�Я�����K���<`=���{���|s�P�Ơquvw�P亠�bM0:�ZF��W!��:�WA��F#�	db�ר���Hmh&��j���烨���ZۻBQ?�71sE��u�B�9J-f��|��B�ο�x��:Y�wSS��:�F���A�'h��/_�K��o~�4[s��w�袋u���y�{�{n�����Һ��k�n}�K_�%�?��?��.Ե�A�-q�]�[�7�0Ft㙔:�&Y��Zv(,���f��m3WKk�ǹ���dM��^�������1:`<�\Ar�����_4J���p�Il��/�oyX/>��>�jHf��g�_�={��-X��yX�>�J�H�&�aa'�h�F��Qo���h��XkD�Aph
Qd���Q�9kbp�bȇo�D�d��L�x
����\μ�k�┲�0�i�?�e3��y�/$�����DD~/Xx��ʸ`�3��[q���t�fX��T�� ��baL��DT[T*Q��3�;1�d"�Ռ){�l8\�)T�c�zU&�՜�C7ȷ5fv/8i��_x�O�{�9��g+�H�r�V�=���?پ�W�IuU�q���->u��l�Ӛ��u�(7�E�*R�] �����_�Y6بB�F�Njo����\��1=��e�}}����-��L�Ĥ솛n������#��Z�Y�3}�}����V+�7�yH;����|�����^mذ�A|W\q�6nڢ�V��	ќ�N������߭�k�����.����*o���Q�t�I��4>^ҷ��-;�~��4������kk���袋t�-�8������蔅���?������'�֖�{�bx�H��Uo,�d�ao�5î18��!͜ܮ|�Q%+�1�SmM��ګ�^��AF2�~�ȇc1��a@���D �Q�Q��[��R0t~H���`H�&g.6Ҥ4ۧ%�m�� Ņ�Q��/�9/Ѩ	x��	����D����t���^�S�U���(�Z
��i a����d� ���
�_���e���p�0
���ld	g��(���i�8Sg�z��E���Y֑��Y�<@A�uOַ��gwq���]�.�7���ӧiʔ�ںu�j�Z��t�m��41���7]�q�0ӿᦛU,��c��!]������>������/��=o�=[�Խ9-u��Ք(+Qs�� �!�~(�P�L�H��°
��ᔕ�F��W4X�i��VA͚��L���.by�&���ok��m�`�e���w٧��\�Rɇ�����'�|Z�z�!����@<*����Abw,���a(Puc��F����ACT� [ f�����uFʥ	�I�Q�D2�ֶ0�1�%Jtol�:�Dw�8Y5G4���ߋ��8���B���r�4f��m� ��E:�:t���ر#ڱc��M����ys�������s���2�2w�=� (O�6M_��c��۶j��}&9s ՟�:�	�DG�0�q�W�̖�8��0�>�<����<���ł.������\�h�V^~��.]���}=[O>��v�ܣ�;O7���4g�%ƹ�?����9a;P`���(j<��-�^����7P�~���J#�F���e?�=k�:Px�ٵ��k�zLE����Ҋ�_�Aw��k���i
�Jp���	\ʉ��'OV���!����RY56wy�%�A!��z�=�aX_�Gw�,��WQww���� #e�j6��4�j #,U�[�E��b:� 4�nF"r/��}����v�55x<τ��/��ETu�P�=4cr�S7��<���w-����?��)T�<����8��	i��y�u�i4Q��}�5�?H6J�&�LL���q���!�9�4����ٌ!r�VZ��u+�Щ��n�>��q��߯�ؐ�Ƈ|��N�����ַ����JF���e����Ӯ�[�a��V�����ӵd�<���Uz~��FT޵r���?�P/�����'�}�������?��}L��v�V��L���#���Yp�P�,_~���M���?��F-���>s�G=U�ӷ�RgW�>��Oi����=����J�Z5�/i��p�N�\')�ɐ c`Ǧ����t��v���tҌI�h���_�k�� +�7�sz<��V7���R�2hf��!g�C�Y �\�*�����:��:h��C#����g[��0����8
D��f�����	�Vq[ݪ$�:�B�] ��� ��j��FnH��L���FL�S[s���b��T^ti�H
+d#��A^�5��������wnA�T��N�L��c�$���+|�,k�niUsC��_x��::u�}���`C�����$�'r^�4i�fL��Ӗ,Ug[��z�Qmڰ�~7X�gt�n�A��K/0��{�u�>�w��)�-kV����nF]B�jY��ՂRՂr��j�v	�N��d]�Fq�D�P"쯠<~*i0/���4Rj���gꚛ>�jC����/�u�~��e�^_O2r��[~��7oz�hE#׭��S�]v���ܡ�[��Z���@қ�*�B%���{2b��gȕ������چ� ����dk�j���X�}�&�]��5&��aS�*F +��f��
�$�0~��X��PA�Ad�#���i�G�UU��Dq �������Q�a �+*�)�7:f�qY`��+�8tdԍ#@��)���!7d��ȵ�g/�k*E��w�d�
���Y�6E�Ur�¨�/�D��ז�ܡ�Ӧ8K����`�F��؉[,����g�u�5e܎�=n��h1�s�k=��Q��a$:��5��}�Bc�U։��� �-����;c+�X��׽�� o�����O�g��駟i����=�
8�z��� ��?����?���o��V<ۨ��	5�t���K-���6I�t���d����u��r�IRvW��ڠ�\�E%&��s�7TDP$#��n���,
��=�b�EtP�����2ܩ�h��pE,J.>�T`�����g1l-*V��:���K.9�o�y�e���b���w�����3/<�ţ}��:y��)󗜬�JU�7n֦�{E���(^*)+���fO&0FY)&�f� �b�TP�!�;�J�:��N�%��<2����ڽg�6n\�����{�>�?�����?�O3�+�����+-C�I6G*.y��n�9׬�J�]���{Z�~�5��]vŕ�����gW�W�ҋ�����=?�G6�!b���w��W�������'���3&]P�(���6m٪�zDm]]��g>�����w��c� y6�TM�f�_�\�u!Mұ�\T�8�)MZ4g��mzC��5wF���Z��
�M�I�e��}�Gj~�Z@4�8|'($-a�19BV�{\Ǹ+ƃig�0�"�P ���1��x��өP����u�h��!ec>���8
�PP�&� �F�f&�����wPwձ��Z�¦_�'��1-C�I��&0-o������H�]�`��5pm�3���h�`m�)� �
�-���c�s?u�b{]��5d2>l�T���fAA��
?���k֌���z�q�sm8D�/+��{���k/� �F�l�]~�i��ѠB�^u����3"�!�G�W'L�Φ�u�[� �(�<��)Z83���P���Z=��k-�c�EdԤ��y��֏��y����k�ж={�a�v�5M�1K]���TE���C�亮O��#�=���c�v/�����g9�&����+��ճ��]���fV2JZQi�{����	�R�V�ַ��(T�1.T���HD�1�D����De`��kq|BgFs�$EJ(]��y}���+
�J���C�����'\�F��{�UU
jYb���1� ��O����dR?#ϝ�	��ˌ5JV[��*U'
�:ꍨ`b<�;j�G����ٮ㉤�O~��ܰ@�ʡ��P������H^��t��1&���+��Ő}�J��5*T���m���:�6��#;� 4�ƜO�w�������Eq?�S4g�,��'?qB���_��^�zz�ij4Z�(�����:�ˤl�|.Ɓ�:��8�hh��dC���S��9M��+�iQ��(-'���kqHd�a�"{	�o���֬��3nFdPd�#�JPhp���!�\9�<O�e��p�|r���. /�]�eBg�lIU�C����.d(^Ţ�"V�*O���ν~�g}���O{��Y��߼�wQ90T�ظ��;�k�����O�W&��ƍڲm�*�F)F��j�J���D��b!ʺn���OJ6JJ��B3����ԑ%7����k��i��;�2ڷ�~p���ml�g>���a�~���t���tB�]{�n��Z=��y8�O�u%�|72��:�x�W^���^=��*�2z�������/��������}w(T��9֬W�����:��e���9m����[��L}�dۻ:�x��fxd\�,Z����9�����U(�	�T6�b�N���¦j����qTJ��Ѫ��m���kJT�5�S�-�z����h~��Z�~Ր9�6��Z.��d�#
���a�C
�X��L�2턻m���D��7Ac&BP���� �C�X 
tt�(������Fa[�?�~�8g�\�}��Љ6��C���g��j���aԘ˵���HI��4\0�$�ĉ�I	�l�)#N�Ŏ,α[��Xp�"�Ց����~�=��c�œj'ri�Z���4�;���N�暴���<~�����گ�C����ao�X�ӁZ�p�Ex�p��~����Ң�Ѽ�����ϮR���ҹS5Z�:�ٚЌ\E�M	��u����B�<��Ji�2S�5�@@�.!֦Mn�Ը�Jh�Pс�a�;�W�ڬ�jV��w�f/<]>�J��ޢ���j��=j똢�._�B9%4.��>���=�}��Uھm���@��	��J�נ��=d����gj�f�&��)d��3<���G�
Ӓ�Oٌ���q��?���O�1�ك+os �R�@��E���6���i Y���#"o����"�)6���Q0X3�d���EϺ�C��}x�߈b�PR�B&�/�=��i�;��Ͱ����'��D�9�����;�z,��.�c��j�P04�&��[��P����Jɑ�7"�y.}WkVw�;#Y7W6�Ą.���皸�7I��9��p���v���EI������.��}�#�/�_�?�s2�w�R<{W��ʒ�G}܈_��nmݹC��}μ=�)����c1�̘�y����q���;0��W�Q�J�Z�g�s�L54u*���_,K������H��/���:Z12L�P-�:��(<��L�#K�_��Z���G�����"���ZV���'��<x]qoX�`�֛s�!��G՘���@��Nj�>kzǃ���Ϝ��+V������)Tk��={>�5�X�����M�ؿ�|��Fct୪ƲJ��A�R���
T@�,�(����<)R�9P�s1���Rq� ���N�W^jF���BG{�t���T۶�׿~����৞�H���'�s�f�7����p���Æ���ޭ�.=O<�~�Ѓ�²8)T�'�޿~G;�m�M7ݬ�+/ׯ~��^~�%�,X������Է��m;y~���q�w��-۶������F�"i�������7�o�]���3.�c�
�k(
jD�\�x���NM�ɸ��j�W��F�7�5cr��[���/��9�-C�8���0oEkc�DB3f�t���l$�����cQA�����ub�ᬒhV�b��,Ry\I�ٸX���_�p ��z�b�תLv�w���M:�9�� ��5I,��-��d�P�i�6��g�d���I�f#�[o�%�Pt3;{:4���CS�v�ޱ56�482jR(�tƤ��3ecH&]`�w!�v������M��>\v�:�����OX5Ft���l��}�g.S��IA���N>i�V\r��>����ሸ�+�u���WW?�XiD3۲�ܜҬ�-_:W�=���9�����5���kԲ�Jy\�ZIq;?G�Rq�x�Q�eT���3<�}GFt�BŔ��U�t)�6I[�RA1>֧�;���w|L�-;G?��^yu���<��^����*���{��K���ˇB�<QS~� �!�B�\��9su����P�����1և8�����L�&�ʣ�j��ܱ��ǖ:Gބ¼9x8D�jj�8Q����:ϙ9P7    IDAT;Y\��	`���0d�n�Twb��3a�h�[}�@��G^�i�(r�w���T���u[�e0��1��zss�Ѱ���t΅���7rͅ[�1�E�BAc�=?�Qq`R2Y5���`�^/)�(����JE{�P�T�9f��3��5rΘ���{h
.��Q�x�0�^��1!#���������|�H�2��ҹg�e���?���zs��G;�+��Ŏ!��*#F�E�/Z��[��G~��z��PS�]|���䢋!�&m۹O�S6׬�����u+��Y�9]���i*���(������>VVWE`م
�.v�F,H�N�V*Fch�����MG�e�a��_��p/�P	�%��w5��J���j�[S�6�L���h͖���}S۲�w�*��g�\���P����o�����#�w�pg,��ʶ=���9�	�8�����@Y�y6�bv�MH���B�A��x�\R6��"�O�l�n�L��Am�@oU����Yg��]{{���]$�p�{�k��3�V�Y�q���v��t��k��7�m�._���gh�ܓ�z�j�y�}擟ԅ�/�֭�֦�/��3�x�\�~�u=��/mt�5���o�L��*�5w�I:��z�������ر�:����G��zz�����:������� ��/~i�����i���m����c�
e%SX�C1ɨ�f䜜q;�[���M)�J��;�G]M)͚֩��F�y�w�<4�7.�#�Y��=���.�t���ӟ���qǶ��}y���y"e�Lz����IP�2���)�	��R��7vzugD�6#,Ҥ��4fH�A4�1F��2�(+%�\y�������/����(|׎���ĸk�z,@�����GqQ��g8)5�J��Ä�G$�*�S *@տ#6Ѯ�nM�:Eݓ�=�Ab��2N"�a1z2A8{B���&�@:RƚY���L*�i��h�g�p	)�\�u�7hճϸP��]�hddX{��I���\G�$���Zq��v0^��&VgJ#�Ԝ��t���PԔ֌�N��(�
�V��c@�c*�T*��Zf�{.�jB
�߱�}Kb��Б����ҡ��Fk:6R����::4��.V�Ȩ�޶M��'��֮���s��s��}xtL��q�>��ɧWٙ�57�WJ�B����vsD(2�M3:�2-���dS>�&y.pY�FUj���eí�uz}�S&S�O���>�����56aUq!�J��\[���C�#�fj-M�.�V��Űr�}9�G@	X?�&��C)��U���}�9z�%{����T�W�偻�ѧ�k���N�~P(b0ݬ#qFp�"7nIч94��(h2�P�%�H�n���h��AOme��*��(�"�v<$�@!����L��(`|2�����;�3�*��D�x.�<RT��'�_� Ht}ސ��S)/>e�HX~��_���H��ho��i<� �Қ�_W�V�y�/��/�}����$Q�
I�] 0-��!���P~�����:2PԞ��J应nhS,�ho1�'��PT��5�9
�Y��6ɌW�՞5/���bP��wI�?xˎ�����s��	"L�|���0�H���J�{��0_Gd"�@|/�_���Ƭ�+N,���bjmNhVwSuJkro��������%˦���VޑBg�RQ/}�O���R5)���
�k���m�4Qn�fP�b�� ͇���Ʀ���GG�]�4d�*����9��8_K��l�!�*���y���HŲ.:U,?�#��Ai����ﳙֹ瞥�]`,�����~�z�im}{�n���\��	PlȽ9>0dE�ھޣ^HW_�R��r��n��*k��Z��y�ع��!ΘW_s�G��]���s~�7^�O<�iSg��k������sϫX�9�0Fq�v�AH����P�dbUe����8��\R�'����Ao�}͝�(6ِS!�q��`�fΜ��o�� ���Ik׼a� ^;v��ȅ$t}���g��F��H��I1X���ա]NB�:� �K��~ԓoyH���j������|F�?��6nܨ��<�_��j�ۛ4::��q��66�O&ԒkV[G�6���'�G��l�1��dk8U5+��&u[�2�w�Ψ
�QI��9�� �N�3:]#)��݈�U�bN���dRW�97NX��;pțETkG���l�C�DZ���ȴ�.��z�+/(��NmL��Қ֙ө���xRV�i��
ypKSֲ�R�C�4Y����۠��6$I�Y	�R��U��4T�z�K��W��H^#մ�祝�{�/�t��5�Ӷ��uݍ7���ē�|Q���Q�i�i����~�E��O��Z�.���A]e���_ؘ��K�,6�ab(
��p�3�C�<C&�@`n�L�S^<o.TPiDȄQ
�2q9�\��j�c,i�"���6�TF��bO�77������s�b�J���
�_u	*�'��g����j�ЧᎠ Aǈ7��ײ��/ ��.N
�o�H �)xp%�N7���V�Sò�c����v~�kR�/�D� �r� x+8�FHK<�sQ�g��j�s��������0W�ɴ��#�B�p�aŜ�߻qc �D�Ooִ������������(���ݚ<cZ�Y�Ҟ]���թ��	��x�ny����Oi��͞`��{<��st��+����i��ۅ� �kS�HIۏ)�:I��]Jf��xN�XZ%�U��N�L���_�s��Dhd�U���0���	�Q��m�B�q���"�RA�v8U��,���:� K�Yk�� O��!��-����1��H��gC��t��5SҔ��D�����J���מ�J,��=y�)T@T6m9��-�ed��Uc�76j�,�M�t�H��y2�:�C���P��`�|�Z��E��044����#�Ր���R�5�[�:;L�B=���a�8�<�.����!V�{z<���T*(��{t0c�,?�Ǐ�z��{����m:�ܥz��5�9Ȏ��9͓�|���*]}�J=��*9|4$&��Yc�8	�tl\�1e�j֤�S�"�0nv;1��J�mU���Q��3��k�ө1�3�f8SU�8��SmBc�G��(M�lR[.����Bf����D~�F�&�O�|�r]y�Z�x�_?�IO�qo��g��u�`��sO�N�0"��P"��@���L�����ܓ��(�͗�G6���7No�	� ��9j�@.�����:22����c�0}P�uhҤ����5��" �Z���
�z��`�u*6�s�~C�Nxol�llH<�
DP��ऒ�@V�u�V� �q��l)6P�q�?��{�&ΆA�¦Ά��!���s���{�|�	5�CҲe���;�����RulH�i�%]U.Y��gj^k\�Miuut��xLȤ[�Q��$��&J �ղQ��Ľw��g}.������Q�$[�-�ڲ70�@�� ΡI�\�᜴���$+��n0�6nrE�����H�QM/{�����y�w<��!��ki���{��������SH��/7?ʵr�*�2e7���:Y�r��&�u�{ ь-;o�������F/[�ѱI��T_�����خ����߇ݻ_�M<@�V�(�ftc�Jy=ɟ�oR���L��s���d`gS�ݸ6Y^�>rUH�j�P�"UfR��4��媒�c$�r��O�ȱubqēI�.s=*dMжjA1�=�A4������̫�͸ZY��yQ�g�� �s��I�&�@`�
J��+R�ȹ��(��H�U`;J<�OGd}獊鼉��8��e��q���Θ��Ԉ�tI�BH��3=�������"����k^�0��yX��M%�,n`��g̙����,�3����MF��\�h������/�F&=���|�b�ݻ�MIlٲ����˗����]�+��|'5�7Q�[�m��W#8=5������5M�̕qy��B����O�f u�>,��"[��gɰ��>��`jjB��%�t}QQ>=�8lm�G�\�R9/��("&�^R��q�u�����U�N7u*�X����U��珢��m���@U�2�����Ag��Ij������|�����ۯ?3�+����)T(O~���9v����mip~I��-���1.�h0�j�dYnj��⭏@(��R�W��'��vf��si���
��I�1U��$�%���"y4�Jͤ19>5K#�>[�	��g6�j�"_
ba,���;���z��C�H��"��)���|��8D"!���x�m7���ǎ�0Y#r&�!o����-�H��'�qA�A��c�1g�tQu6JY[�١�>�܉�4�z��i7g�$�Ջh���������=mHF|8x`�� d��=�!0�Ը��C�;78�OΝ�׆L����L�ŋ����"X:��"&b`�&\Ly|�����e�̳U@9�$oNC\��f���9�rR*����&��a[N6��+�[ݯ���\�*\)W&�d��ۇy��kl�.U��7q,PD�d�-��~�B�"�(}9H�q�t�ю�&YdF��\hj!�5����܆r� F�6�����F���E��7	r��1k��	�#)G�~ �H25Gi,�efgx^R����~�zm��+_�:J�<XԞ�¤�;��򸐈��f�mԄ�p���Fo��2+�=��Kr�B��t��*�Չ�Ldpe<�Kc3"V<D�۰q�VL�f����h���5k�bժkT���}:�7y�;�c'On��JC���d�cfe�FD�v�9�N�	ω΅��1�X��$ͨ�^��pp�E��&Gu�"n<|�o�T{��.\�~rE�b��Ϣ��F(�@�9)��?���ee��P����f<c����9ƅ�+��бb#�%���&�
A�{)�>R�T4z1�MQ�Wn`up}"�@�⼞M�%�j�C�0�����"�2�3��G�4���爸�I��:@�O�"�?�W��exIXgW��0��$r��r'���X~AżI�D��g�_gD́cu�����he�r����ZTV���ma6ܚ�T p��t��~�����x��-H^e1��ى��cx�c�� ������$T�{\:���s�
'�G��U�?�A8ى@$���A�!*���|P"�I��АS�CSq��5E5�g�.�V��Da��!_@(䑒���.D�$��I�SȌ`j|HQ'$���&����f�#!��Gu�S�[�4���b*���2E]��Y�D���%�hMx�	Tp������?��{���s�j�)T�4��ϟ��Ѿ˟��|-Y"&LD&ԧ����Ɂ	�ٹ1�0����́)Id�0m�k&�.�*u¦�P7�>��"�Xs��s��	��(J��,~�􌒜����;1�	���� ����a���xv�1��ɮ���ɳLi޶y+�mي�/�烱æ�jC0���$R3َ�.Ad�J�0s(e�ډ�i.�f���(��Ɛ�y�$ɾ�	�d�G�D�v]8�d�#�U[2�ӧ���)&'�А�>�C5��VE���%�"O�.]6Ax�P�P��u��Q0�-T�`5�p
�'1=�l��Q-���;��Y	&V���N��%���q�uY��s�b��p1&ɒ�y��<e��7<��̛F��QdT ���{�(�H���[4¼!�	׵!������5���B�`�xB�r��p�R[�
f����,�fE:e%;��'�b`�߄���*�w��\��ia'�l�Th�#�`q/[�B�C�N��8�_B�|=�,i���5����!�n�LDB
���4&	֤S	�L�l�
b:�RYx�r}.O���4&f�@ ��;��|��l�q����8����Nc&�q��pL�b����,�tv2G*�
��$�53Yh�MJ׈��q��՛�^��؜��:1ɳJ"]��ሮn`֙���*��
�P�h�OZr�*6*MI�3�6���(�{,V����a�j�!QB2�o�"�e�|(���V� ����f���k�v�R3
�F��ݼ��o*f���c<�Zso%S(��G��b��Q'�ߌ�,7D�5g�U�&iޛFxv�5(���3��]Z��g��BE$T~G,��@�h�&���������+e�����~��Y���"��;,�8����"����#_��38ׯ�h�B9�.Z� c#�����ҕAD���׸p0���n���[������W�3���N�"M�Gj��x_满��ׯ���*Ą�m����f\D:�2i�t:"��a������(R�]xx�4F,�����L"�I�:���4;�����m���]�xk7����&	ary*�ȵ2|�'�J�5$�L̎��9�X�c�>�b��S�7\��swoX��;��NG[>�����o�P��hw?w�g/�~�X�6�|��.�G����qu�~�(�R�"���bI�t>$AeEN�t��08�t���!���y,�"���n+t�0���X�ĩ���f�i)[�0��
�qA��:Z�;�}}��F���J&u�s� F�1m��L^��ꮙM�	�pS3����#!?�$�u.�<3�t��Q���x��v~~n|�Xy�h���nF����:�>"�*&�����9�C2�ǥhkk�qP�Q�ǜC����D2Ǎ�q��	��a�G�G]V��"�7h��s�����K�7;b.�����V���w.Q�vo4 cAd�-�N�7[�8$/>�? -q!V�-�t��.�Z�:d9?�2��(H	�hs�'�;�!�],޸0�c0��f&��"�p4&��>�0-�i�D^L:4�k򇂴��2Zu����[�zAo���q�~�E������sgV��{�Rv!�����*3xm���#���#���O
��
��h a/�!$����)@�]7N�As�y?.��WF�2r5jW�c*��d���LI���b�Pv�H���>Mm�<<��Tʤ�����[�����{��PƓόx؆�A3�r�E,Β&�M��KgT ��!U�Tk�G�^��ΚE(��]<%��j]c�Y~�CN5��1-��uI#MW]2�<���FC�ʬl�k�$�Pa�o�����&�����f�!�;&:��BC2�i?����t0=�
��8�)Ɲ���pQs�,u��ZCΓ&=��3*R���u������h^���|N�1�i�,�9Rs\�������lQd�4�d����+�8*1���%q��v����wɬU$�2���UxFu��2�H
������!�X�4l��{�1WD8�@$F>RV��ؼnݼY�uj:��}ǚ��_Ma��C�m�����Tgv-#x�{O�*'囍��L�x�ё�����|:v6�T:��\�=��x���R~��b��4Ο=�Qe��A�D�8��zG�(����2o1._�XS7�(�e�G�5E^b��A��E�SGK$��� :Z���Ɍ�؉=�:x~���������&��Ź<�'�g�w���y���'?��כst3�R B���D:�?�z�o��?$W�͛�n���3��S�Q�n�*�_.�$@�z�E֨��f�nl�IdB�+/'rx�	���
T��4�c +^��B����ivŠ���}�<�ªTV�G��l�"]�T�m`�x4�l�fV�cC�d4�$\�j���<�Ͱ�'a�P�!@���&�w8]�^���Z*%9���S�[/"t�����
G?\��ϝ��?��ܹ�p�zz����g�g%���ɓ�Ig�Y�<yZ<x���|J�J+Uu<;?W��@��7v%�ti�f;�d�b.�<.*|}+56]�����~�)�9�� =�2���]�B��t��݉��a�����z�y��ϝ0P=ϟc.��I䋟3$���s��@j�IVn�}���"@3ԭ5٦N�DT.q�N��{���	�����R�4�F��3gN�&��ڬ��k�ΉCp�EֽAU�Us����ԣ�c�B�8W�X؃�A    IDAT��$�UG�^B��A)?O������1�[i۔�+�E4��U��8@0�z�VE*�Cz&/�o(�h��;�b�I�A��L��?�ŗ(J�����K���o7��5��c!j�{C�v�����to"vv��3}��y�,0�;ǨBT��gM�8-$�P	W�Bi��|	�t�y��g��j:��i�Ǎ�&tW�0O3�!7��
�Qn�����FGD��tV�꺲��H�k9��./�j5�C��r	��4B���ذ�Z(2�Z���4LE�b����c	���2��Fd�ZcP)�Zu>M��T(�b��b�%��b2rJ�9i��]�cq`�+S`a�/ei�v��L�Q�QgUk�?@_.S|h��D�BT��[�z&Ë��U0n��8~�U6�����ܨU����r�8^WS��؈�d�H��9i��Kc;�U�ݲ�7݄r����i�8=�Dk���)�V��/@8ނJÏ�L=�T���r�U|�u9�V]�&5�G[K���e��"�ǃ:�f9��#�+����";5�ɑ�pU�ضy�����w1p�<ܞ0FF'�7i�b���,m�)d�ѧ��^�,^��E�Q�D�)�Q�)�Y���Fh�xђ��)���N�<�Tf$S̤_\�bɧ�������F�F���Kg>�y���3�bÍ,=6(ӌ�0�����T$,���y/o��lGkr	d�ˍ��WJ�2�aKE�lt�$˸9B6=�F����z11���v06�����.NV��՞��`b�]��%y�3m$���u����2�Z���@�Ft��������@�e�ۧM��ߥ˃BC$[u��B1��]�<T4��M�C�
A�^�\�یT*p��C)�4�C(�Gu���-��䉣&������/4�X{�*���?/n���P.UT�d	�9��=�C�C��%]*;�D��[��1��N��iA�9C�w+=&j���C���ۍ��n%>�|��,B��7�X�bV�\*5"E�]�z<����g����Æ��d�pS�q�����Pa�h���y�FY���s.Z����#D�<��� 3E�_���%���M���<&)�
9| Ǐ�ڍ])G�De�j\� @�ܹ���瀝���]�a��94�q�B��OS�BV�ϨPa�&��m H�z�0����9���v3�2�*,���+�$.��p4F�m�S錺�\>��M��AU�Tԯ1&���,��Ȱ�b�ȃy>����ܿ���_����R5m�,dy��<��?�.�Oca���q�&��	��;�qk�6�qtY�&ɲP���^AŒ	��b�H��a��-��r����󺲄ZkOO3�{D6{^&��1
D�r�T�9PQCYvwk���,��<95*^��r�,th4���\��x�<7N��������kL�^��P�R���f=d�!Y�䋔��� ,
X츌3-�+�ty�JL��DYorc�tl8i� �X)�\F	��yb����b�����-�˦D�[T~I9i8*k95n�6q]�<�^�L�u�(ɸ_��*�e�F�t�u
^�^�:"� �|�"��U�M�̹�H�u���h��(�����y��J��}%)� �=�B�KC���4"���Sr<&y��r�%>㩊����R�4�S�L�\B{Ko��ͺ�	���0:6��键-�K^�|�d32n���X����,�'Ԇl��R�*ɒ���7��h
y��FK[��:���2�����,�؏�������x��
��_<򉁫�?�E[[c*_���4<�(�RT�d#7��Q�b$}�R��>�c܀�\�n�ܔ/{%d����h0�baa�\k�[�;�nǋϽ�c�O�x�����^#qe�z0E���t&��W}>��k~+{hF��U9S=�n��(	�)R�v�j��ȉ73M�Z�Z����V6�/jT�vI�ϴ���4�!����̏�A^,��g1BCt��Sk�dH�4L'C��h�W9���et�Ĥ���n�����������"pc���җ���-;R�[�!���СC��׾!���<~-����|�n��2�Ԧ@�PB6�A>W��x��"��K]|'�Ԥ�Ɯ��أ�>K�����ц��Ǚ=�)�2��-_��+����	Η����G���~�A��NN�u�&�`A��["�S0���7�Z$�-N���NON"ObͪuX�u�C!J��2NݫQ�{dc�Q��?%�4�;��0�51>��}�gaKΏ�M��9�C`�x�Z��kBy����B�`P}�q���B~Z�{�w ��V�����#E�	��&5��e��8�Qx(I�~uV%�������nT�xBA�)ӥ{��'\h��7�hĸ�V�F9b6CS��E��=K&���C�w�$��#�*�\�I>�:G��T#U6# �1ӹ:�ܤ�~tbB�I�,�H�e��^QRs� /,�1��o:_y�j@�V#5&B�z�Q��K���X�d��̟̽!W��gl�����Ǣ�)���A]Lgq�V�mT��܄�DM�(�Ϟ��(�R�Xĉ�?��a^�zjhtk�O��N~�D��N�C&^�r����xS�N�ȣ���*�>��6��%jR�i�͑�b�?���*�`��ɗ�\��Y��Eveк�$��s�#1���l^�+�[��j]Ra^s|(	�TQc�F�fy�h|6&�Td^�BX�{���%��dy��Aa�-۷c˶��\���K#H�u�Tw��p94!��+�7�R����y�}�?7G9<�x����H4���>�Ͳ�f�,�P�o���KzQH�����XܓD2�����h��E���޻�����142%�׹���/Ž�ԩX��W� �pwT����oA���0�� [��C���jM>Z!t�'�`��¡�{0==�5��5+�}����������3�cz�K/��t����+׷x"^\/��� �3�8{�I��Y���BM�^-�Y��z��WE��nI�d>3�:gb7|nF�Wp��;pכ�������z���DX>!�}��&O������Y4�e*�;6��*�
��N�K�9�r��0��.�D_�h5��1c��[m-m��<��P陔HO
�#2��I��?z@��?�����t5�yn��pC7���10���([�⮻b�1���@8?3���0"�:z:�q��9�tX�Yx��+V.�W������(������c���W���g�g�x�892Ae�h1���;,�B9���A���X��mq�4݂a�[�;��"IZt)StF����z�6'�X��+W.G�)&D�P��D��ׯ|?{�	�ON� �qo��H����UQm��@�[��X3��2�Ɂ9\�jV-_��#�E��D<���������gZ��Ǚt
��^{uN�<.8���"��3	�$��eR��kpq�9;�X�$b�Y����R�t,޹1=��YD�O�ܙ�d�����`G�N�͢���O�I��[�wHwZ�w��C�ɮ��C~7��"����hQ�57��k>�aJ�)�Θq*�&ѻ9j=3���G��.9�a��0������/�H᫩�qyonEgW��Qt`�� ���Ѳ!!�B�?M2to��t��]	�f����*52��V�
�֢1,�㑸��Y3���J�vr�x�y؈8�j,�laO�W:\.���� �(�-�����\�i�B�[g�7��M���nֵT�E(�w�ʠ��E�	#�H0�hJ��QPYʏE<�Z,0�j��}�W��g�6�ڑެd�h"�1�Y�󚬘RGMn�������K��`X�7\*�dG@bz�(�O$��"��-��*�H�8��y�;,��:��$��ˉ�%��9���w�n�&i�q\�B(тT��Kc9����6��J(p�����L�IMv�k��ޔT���ro�p��
�+B�����hO�p��L^�����h�4�M� �籖�ۻ@�T*���.�RY`q�z��)�-[��X�~�G�p5��45?����U��
7��.��A$�5����%FwGw�Ӄ8vt2�1xj�s�/��_>�?]���KX��*�F���S�ǚ>�9��� N�����?�;�D���d�_����'�!<���9�&��/���dv.�E��X���2zkkM���@!���[�����`דG����u�h�i��yW�A�d����/B)7R&yr���Q�BEF�h�Rav��ZGU^��D�eퟌk!�1�-����/�i(��7���{�WR.Q%�.La~���.,l�p�`�q�:"�8�L���r��-�Ӆ5�F���E,:���Ep��!�q��BMD��5��}�����;&r�잽���׾�Y�� �f+=O���k�%՚�u�27]���Ϯ�h�\�@(�ǻ�A7���l�=��N�n9��{`"U�6xl��'���aނ�*4���/�]���+5�c�MN?��G��(��A:((��:`�S��f�Q	chh��]���狜�k�hUk[3�(J4R����g�c�"E�>}
��s�����E^� ;�,��q��)�ͦ�ʠJ�x�`Q5��zSi#,U09��ZG$�y�^���ϨJ�ǌe�ŏg����л,�i'�����
��]��C�7�a;KExG�@5rF�E��1�$�ͭR���E�27a�=+��k
n�D�4���b~(-+w��渕m3]��F_,�X��w�`^�|*.]�(����Da�~E)�LKLru�1L��N�T����G6�|�s�#�7͒�L���+ɕ٠��8���u��O�]��p�H�ymd��!��xtL���eі�`���q��a��;i��(i
K��&����\
&R�1��>��� �%C_��h|+�I�i��f�Ff��{�/����*x��
t�����|֟I�&�?�X�T���2oL�%�˪�$�q�~)�.ttu��hJ��A�l~�ёj,`��|� ��Y(�ѬC��g��i��X���(�� ����;q��[�J�h�04�F����$��k]�p��`\���?J߅�Q*Ja��H#0�h�
EB�(r��&�5e�c���jh�0z�4.�F�U��mX�b>��	h�������
�Q*���ѩu��sc���hn�P;n��<�,��;���8�5/��.�X����
�pq�A�=@S�'���B�:��G�w�KBT<���u������߹���H1���o�P!�23����Ogk�VV��Rx��_ �&L�j�U�tǙ?��gg�®�SK�\p�UwA'�Q�!����hmI`ͺX{�r�l3����?�/���<��������\��˖����*�<0���W14�ɏ���2�����ẵ������K�h~/�lڟq7-Z$���|�x�e�߻M��x$��oĚ5kTMOOc��%�YqSZ�l9�z�}B3�ǧ�Q*�������chiiÒ�K�r�*,Z�XP��Gp��1�"� ht�ẍ�t�ds�߀pȇW~�Nڇ��A4�}h�G�E����t{䃐��5���/Y���# [�J{���W����ް�����Ba�z-|��؎j�w��vq��&����N����ؑ_Ϫ������bŠK\(�K��/��ŋ�c��5himBOO����VJu�/|	O=�K$G�5[�.?���*�?��7�\7J.|���ϛ�c߷�5���lzɢ�����u��+���ẅ́@:�1��s#����ѣ��aMA�K$���r|����Ą
�
ɝ
D2i�aq�����A�7_�נGqa6��o���x.�hS�DBc%J��Aũ!D9)m�i��p�L�s8j5�=��+FA�ߤ����i��O���Iõ��tS&��fBq�l�� @'���dg�q%�1�Y��	��-r3<�����5�9;p^��!O����Lr��`�I#��Ajx���4����@$�h"�l��elv�5���.f������<�{����h�$�Tʑs����6�	TK����т�=��xq �.(Hj)�I����T�p'wF!�.�8\W�^5�{�hY"8�K*\����Ō�X���pm4.�91�Y��Q��;2ל�X�H��-����ؐw���h~:���cb��k��	�4Y^�4��*%4'�MfP��b�F���`Ǔd�gK��x:,�M2��_�ў�5Q�Ӡ���,v�ts4�d5�gj�a����n�m;oQ�����'fP�q��%Nm[����"�s�c�˴� nQ��]�"5~U.��Q��!�t�`뎝�5�����
�>?����|�N�{�����Q���5�����:���6�e�.x<�K�"غ�F�~�y��y+�����_�w�;r���'硩k=��x�X���1�eq]Fw2����ޖ�1?.\�����PʡRN�[�����?�fM{�?*Rt/�:O��>��h�O������2�B粵�b���Ϟ{y��5T�a�ı/.^�X���o�,��Q3�/�K~
� ;�:nޱ�V/�<g��hND�U�}�e���,� n�m'��ج.�S0Qѳ�� ^=p\U)7�X4$8��ٓX�t	���C:EEO>�&:�cxx�tt��Q�D�
���C����'t�v�m�'�N�s.�=��8|����������%=�BjjJ1�{_݋��!%tr���Nahx=]���Չ�{���H���]�?z�C�LϤd<�F/����g����x������g�*��ݞ%��H\�d���/`Æ�$������P���'��#�`
r����e)]Pv^�,��9�}�\dDp��6�����l؜�_y�E\Tq�����,^� ��I����b���Z ������T I��b\��X�/�5�'�Cc-c�K4��󹢬���^�4������k�]��a�����"BT��y����Nٜ�tT[���� �̗�NO�=�ED��'0�q?�3��y�J�� S���e�g�ݳȠi�6r=�*��}4�(�HRh�ϳJ��Z���Ľ����XL�-F����BԌ������̌�9�Q��%����'�iX�u�ƞ�!�~r��=#�@��>����?�X�/,��5d+�T�nmnW�ʑ���K(r쪻�����B��;���'�u�p��*7U�9��k�F��J�� �}�^�P1�mrT�y[\Ru�a�Ҧ^��-*��4��{�ޡ΀F��-qdS��AK"��yzjQL�lNXH�3��y?\�n=�}�[t��0�����!�'��!=���X�Ԣ(V�nϹ>��&��p8E�#"��y�nϧ�Fr�BX��:G�wƜ�h�6K��y�W�������˘�0�a�K�8;*>�1�u��MNc�I��4k����~�ɑ,���#e�8���cB5�l�p�XȳX3�h"]*n��*�]㗠ߍ[w��Λwh��Le04�F>*#�*B���ڻ� y4�V�3u�ZI���8����ۖ˧�T����a�����`9�\��tE��A���.L\>��'���ƒΤ��H�eBy;���F��^�feC?}F��{�_�\'�:�#�u�[����������$�e/���b�u�1�j��L�#֪
��P�>����r��@�BSթ�k6�������vӲe3�N}�*TB��]���c�>oj�Y�i3N]����'҆��&g�
�b���fU���Q*+�\�"I�b��謹��@gS��w���Su���gqi��悷�7�x}d7^��6n�o��v�3���c�� "�$֬؀�t�Sg�#ǅ&o�3�������v.���c�<"8�����G��Ů]���/ �˪�x�{ނ�?�ܷK�.�MEX�ɧwɯ����;vb�u�����Ϣ{^>��O*��GU�2j.�X��|�;u^���o���>ս�=��5+��[��v=��l߁���wcrr
{����)h��";>���.U�
)e����e��ï���+��_>0�d\99��R�Ё�����C:\4��[�0��Z���X�U�X��nW��    IDATR8J�yY��l.&~����8�
�Ю�~��t�&F��v�F�@�"�����b�84<���b̺[���Z1�j ������k׮|�ל�����ի��ك���]� s5,��|+�/.GgV��k�t����&u���E9vT�iB�*��\���(9*�=������B�P�A�\��1Esf�(�0�"8;�?�!l���w>>>�b���߿Q�P�Dt����o��d�Ų9&n"Dx�����{����P����Z���4�s���3Bn�Fj<n�_�%��ȱ�yb����k]�0���li|�D�/Vc442�B��b��\���|�$k�[Ă��{H���nm�DXH	Q�����AT
E��u^'Kh�$WBI��� ��9Ou
W�#�B^�,�� ����U�\�f��g�p�� �� z��d�@9:e�����|�?#2��+���������(J������c��,6&D��#S@ِ?nؒ��<9�8p�`�7�p��f"�:�_�GS�Y�9��s��Q���y�Pb���\���;����Ǚ3g4V�"����	�7�
)?����=~\�"CA��L&�:Gy� r�.a&�d�&.C\\��5*uF��-)���fl���;�;A�`kU�QY�lߺ�AT�BT��1��#ԶL�J Jo�MM�&�Q,��ù���<-Gj�DB��z�h�lܼ�Ep�� �9����Б���0>p�-~t%�y���锰�u4���N�@�7�y���>����w��N�_��zZ�=���x#�Ƨp��)�L�+5-Ĳ57�PMgQ�*�t�}���g/^Ɓc�Dޮ����.H|����t��%��Z����ɽG>����]�t�������!�|�a�|	̔�t�
O ����P��|�*��tO%
A� D@��O-��<��2��)t5G��Ƶع}%v�>�^x^W�lFi�o�c~��Kػ�0n��vܰy%v=����%2��n_�p$�B�&T�B�Q%'���S�҅pϛ��G��3�<���$�w���hJ��[���|Fh��t�|��ĳ���<�M7݀��?^}�U<��.�~&Ƨ0�B������=��(_蓟���ߏ��{��H*۾c��~<��cx�ɧ�2��ƛ6�|/��2�����ƽ�����s�=�y4=<�j�<�<<�"ڛb�6�8�ק %�&P�ښ����&��♌�����܎H8���}H�$�P*�B�����EG^RҘnX��ȑ�Lg:[C���6M��M�Ջ�5,T��I�h6y�	*�If�k��X1a[��\B�d�;V�\���oL��I..���!���EK��KMM�X���r�ͷ�w���$��G������C*g�Ôf�3[�5����F'��w�����#'�G� �O������Xr!G6vs��\�)a�&Í�rR=T*�p�!u���t���c�̞=_�n�T��?��!�,T��4�q�!Ds��C(��av�|���U��XL�"�x��q[�.Q2~W�2�@��$����ō�N��>�ul�&��-�Y$��1�_\o&gR�=R��IG�D>��^�\�ԉ�~��!���#ې�IC�f�Ǒ$K�F&j�Z��O���ߩ��R���Fϑ8�v���^P�����K���1>|G���0�[���B���YyTUZ���p��#�Mڼm;��o�Z����O��ӧO��"��R�%��ԬX�479�>t�8��������y�����9�
!K���=�aYas`Ta�¢����6lAϟ� �(���h�O"�mvH�'[Ԁ�}�M�|����wC f!����"�6Ȓ�&R�I��!�X���АG�s�v��p:��`d2�t���+�H�}�.EӼ�D[����� 95�)�9���ǻ��Wɘօ��˰�7"�܉��������B{"����@q�"��~,�Jb����d� G�?���4[�|�(.\����$��0<xE�jI�7���i�_���4�e7��6,^�A��3�X�4*h�x��@[����.\���GQmTQ��G�-��/>��/m_�������CTN]~�t��Yo8���ێ��wi'�b4�G����t�pR�l�Z,�2͓7ɬ\,#��9%B�g�q�-wފ5+��³�b�="�ۺ���ؾ����^���5��DKG��C8q�<���AO�Q�D����P+�^�#tcú����Ç�Įg�B�T�|���ݏE����_�������ۅ?�_02:�o��q뭷��;ވ��~O�z-m�HMϨ���O��^ƿ~�KX�p1>��b�s/�����.>���x��x�{߁���
�$Ɏ�+W���c8��/�嚵���?�C�����G?z���(��pч!=���=���Pnv�1���ĩӗ�F��.`����9ɑI��rXM&[��'188��V�m��j�y)�t<M���M����-Hlb�3�u��\�^���2w44����Y�F���NOb:�N�����2?+Isr5^~ֹ��M��2�wP煅.�e�V���aF-F���YZf��� D�\���h����~�0GE�mZɇ�D�ZD	�J��}��abj��(��D�Z���!A���<{��x��ư*�tS��#�C��,��XX�s�wm�,�	�;}ERXu�P����7����B����G2�Q�������9���ѫ��,%��7��p��a�LBU(I�E�1�L������D���uicq��a�g�!D�I�q��L:���⦟��#?"��c�l^
Hd ��>3��N��rsX9QZB8��XD%�{r�4E5G�arT<�+ꜙ4\�-�:_��i�����ʆkV�M�l������˘�E;�T����Z���,A�jI֐�6ɱ{�oǻ��n<����k{0x��?
/�y��p�cV� �&%��n(g���NU�!�h3�	���b$~�����kYƊ0�!ߛ����g�{�{U����5DE����E4��1�4���v2�E���E�o��Ui��CI��Hެ\ʠ@������Dh�	�5&$"�hm���nڄM7ܨ�il*���,�U\��L-�h�
$;�I�R��H������0~��%�˄���SQ�Գ�o�UW�"Ԗ���υ����{~e
1w��[���lD�ٓڷ�Z��b�
=~#c㺾Y�w�̓��=��h!�Vo��7�����8F'�8y�\�P+��ـ�W�P�$��F��r��38t�S��F�/j����������}����v�B�2<:~N�<�:��(�2��Hb��+��ꆂ	m�$����i�p��ηݎ7��g�����\y�ML�}^x����=���{�z�*|����k"K�Pd����A�)t5+���B%⚕�p�����+/�g�U�������q�����?+�تK��G���}�ض�����s/�?}�Q���B�����1<�կb^�|���> �?|X]-��;o����[�����m�v���~G�ŏ~�#�X�
w�{?N���w��]����_Lq��f&v7�.�����Ø�I��@���B�0���5Skk� N*1X�����*��6�<a��ڢ²�e�� (|O�������E�6cg��E������:vG9�<����#m��3B�a��Lh����hp9���ܐy,���mH���82�����땢L�7D.ʩIr�"���Mظq�:VA�!SY^?�%2x�<,^W�޹��Pi�aD��ղ`!W�0�5�R1�FFG���8����R� E�Y�$ܒ���|-��2BƼ�����)|�
S�s�10(���5�h9R�s�)�L�!yip�h|�$�wFs�N��$vR5�ɺ�0|���N�9�P&�H��H�Y3���ު���u,�FN93��7��8z&�r��*���Оר�*�E��"��w	�)F�k���)׈j��y��k1n#2�g�C���I*�%�L�
��x�����!:�H�~�f3궉��۰����͸|���*��^B<DWw��g\7���>,0�5��UL��?Mݭ��Ac��N��Oq��]b�h)5։O�F��_|C6Ϸ)�v���e�C����	
"(D���l�o,T���6<־ &��h����3i}�S��X����witm�A!��!�~��i�û�q�����;�\s\?T�x�'���]X�t�qc��i�F�p�"���T�L�+�"� Ҿ��%p�I�C���[�c��Y��̌gE�d�b���-�<4)28|��QƧ�38s��s��n�c��V������(�e%�G1�J#5�S| �zƫ��7��Gc����H�8r�}��19�G��Q���uU�k.d�g�i�-���֠
ϟW��Z�]������}��mD����ӿ������]����:���K{N��x�|L5��[:c���G笕鎬�J��6�;�����X��F(+`��u�����cx���%����~��q���Џ^�S����o���m^����'?A��B�PE2ىR��b�vNn���b~�ei�7\{����x�=x��t���=o��5����_���'���ތO}�ؿ�5<����Չ�����z~�����f�[6o�Ν;��K����==���|B	����%��"���w��]�K~��_�JIoD�v=�y��.\��}����������2�$�6�r�u�����X��	T
8v��3(|��
���Y���f9~�t��	�uvti�`���T�CB�).�\�nV�����Xgn��.ls����}�-��&<�H��Yr);E�.:Ez<H�'�Ϧ��U�w��<�+�� v|p���g$�EuSR�0K�^ט�����Y'
Ơ+5i"�߰Q���xU��Άr��t`m*쾹��:Ap$:�(�011�ݯ���ȧ�}�z�B|��x>d�%��'�[A��h(�.�33)m�<f���L����2v�Rfn&,V�d5�n)W��S*�&ȑ�:��;
"B���'�4�s���7��YT���d�����/�/��9\)+c����u)G����O6�1:<���A#}#��Lí@�"����N�B�J��y��֨A�����"���λq�7|�D����2,~=�Q'<"���ê��
�ш
�<�L�&b�M�N��܌�o�u�K_�z9�]���p��)����m���EZ*��u�{�	 d��=��d�]�N��<�0&�&����07~�H]�����_9s���e{����]��4�
^g48��:�n�@;JD��2�Lf,g[[��w5��R�F�R\!��-y6�c���MyΠ�̯1q(~��Pݨl�i�#2�'Ë�;��r�	�N�D(���BE���Ru�Qٸ~=6�x�F���'0�*b:_�h��|#�P�R$:�!���2�x1�<� �(�J�	\�ЇJ%'����x	���m=K�7`�3*�QC,膻4��G^E-3��۰l~&G(�bɒE�OX�
u��e\Åt=��`NQjj;�m���q��q�2y�N���d�U�r54�q����_��r�2M߼h��0/D�z������VK�#k�7}���o��*�^_<��;�:�?��/Y���u����w�Z�)�<5��L���1��ef�T%��O?V��BM�f*<`w�n�t����y�"��W�$�Y����$C}��]x����׃<�A�~��g�SY�./_�}}����}��(�L�B���
X��U��mÞW��&��{����{$q~�k_�ї��N|����K�=���v�{�]���kq���Ν��u���Z��r��a,�]����T/�~�c��9�����m۷��_VqK&�|�2���ܴn����?���'��?����DE���B�����64�yͱ5�uL�[��,�=H�7j���i�#�4%�Uiy(;f��xɏ�3�e�\dn�b;�]��MG��v�s�3wDd>v�����w���<���g&ħ���ұs4��s25�ZR�^�� +s,�pk��ꇏ�d���,2��e�k��}����Y�Z\g�!�јb��J��ј|q��[����E�o�]�4�{����ذ�0�
-�Q���.�525�Y��|��*�(1��-ܐx,��w���3��j�"���))<8�'q�]n6KT�%�N��4Fc�k
!
�*�rl�?�����̕��.��(�|'�j��?��h���L��-��4�uU�Gv��Lp^,B4,�M7^������/{�|�[�R�3o!�Ʀ�	�Q,��>e$�����A�7�+�!Z� �ś����,Dt��Ġ�03S�y��ֱ5orH�F�D��)W��T��,��:�l�*l*��֬X���gOŉ#G0:2("}WW�<��j�23���I ���7�	�6mR�b�-���?vR�-x�Y�ZDS7^��I�ef)q�ci�E��*�8-GĮ	�H5��j2�=��ȑ�
�N�81)Ն�fUj��P��S��9��)ɘǷt�"!E\S��O<�����������=�+���� �]F9C� aM"�J�n
!#�����ĸ�("�v��L��������U�pӦM�/_�:��T�0>SD�D�u�]� OH�?A��)=/)3����z��7�g����E��ŘH�pe�Yh�Ǡܰ!�wxF�b�u�q�w����F{G��)��O_��]x��t�C	5Nc�A[[ʕ:.�"]�����y
^�5uc��M�\�3t�.�w,��p�I�clr�*TN�=��Z)=��7���������3��=r���❽+�X��"N����L�
��xQs�i��詺��H�#��պ�!Ѩ�!�vD"nsSp�Jع�&�_��.29�J���x���u��x㵸i�&,XЅb�ϣ���+{�_Teͼ�D<�0'~�˖`��k�w�4~�W1�t� �n�Y���?{ǎC8�â=��M�cd�
�;�E���M7݄%˖�:�RF��k{%��U��p���s��h��R�B��W^yI]���~�8\���ט��;\�)�����q��a���*J��|i�|��YĽ^�7E5�<|`�� �d�2���L�*�FiËx˖�Z�x�twϓ�=�Aɏ���ūq�sQ�?�4�<k;�_^�����:G�l7�_-jL��eD�������V��R(�PK�>v9N<z��N�~	�����L�iGY�s����xGk���K.��n�5k��}�z�M�T(���,��]p1��ԒA��!��6�n-���R���sODeȈ�{����gO���~����/���Q�N�q�y�G��x�Ft�n��j���������Gq��9��M���~ �2��Q�@��r��0�ʞ[[\J^[2пq�\�(�����$��I�n�T��葈�ݜLc��U���|5)�:WU��wk[�6//������߄���_�*��_����/k�^�|5N��c�X�`��E�P�Fe���1���8�T��m�x4��&�}�m�h�D\�t�K��!ќ G�|�k�Qc,A�� |p����Xr6�C�l�P�jk��ބj1��c�|b� �vI�Â��
�;�m۶�C�_�e�f��`8k�"��q�)!<��c�ʠ�7v�y�92l�֘�������%�
�u��xXҽ]ر�~q�O�Yȟ��m�w��ڵ��9�yfi��Ȃ�曷kD����j �
��x����BX�Q�+�@M���bb��M����p��,bb� Ç"������1�=ݲ���N	Q!ߥJ�PЄy��X�d	n���!��2�r=�+�id�@՗D�}	�m�������E�7�hke����EE�pd�.a�h�	ɦ6��b�D��$w��Ga%���}�pj?z[ø�����p��1D�A)����E/����j�Y�P�l�b$�)ǘ�w�� ҥ:�9��1�?�p��\�	��.Lg�(R5��=�AG���R�OÕ����ң�+��_����    IDAT��������Nٵ�������o����>}��rϪ��Ŋ}'	��"����S�0�5}�E����20x�0l���d�s.[��
{1�N����6tu�jQ�M�,�u�Rڰ�����=!s6��3�JE>���<=[
Z��[[��rtBnL �x�Ԕ$��&����	�peh�H�j�����[#;##�33vvq�d'DOhutt\7*_�].;�$;�hTsu˴���R�����=+d��L6KF����]+��a@1��ϭB%�w���c�^�r1�!-�xtr�\3SE�~�u���3��ۻH���a����ߎol�b"m���������7����!?6�F��A[�~l��L�n,���Vdh�ͦT +����fn]3�	*)L�JO*��N�q�,W���)������[����-��z�N�9�"���,V�e����,��X�$���'7":�z]?O�_����������(^ۿW�x2f84$�V�8���HΞ��xHLe�F}�z����b���o�����s}6�M�OMI����W%�,�blbR���
��YdU�D0#�]Z��;|XB5��aW�".:�_�ʤ�����Y����8ۂ�v�DR�r#��h�"��̤7��V|���������6����Y�ߪ�kq��y*<&�������r�%�_r��6�F"D���j\ɑB����*)"1��2���"� �܃����9����)����e8�BZȝ��*,|n,hoA2����&FДK�<99���I]#"��C;�c�-�7K|�����8�,�F��>��.)̮I����Θ��q�c�U�&k�P�����>/f�c
�g�[N���C���B�W����-r��H���v뭷h�z�
5DTx�B���p��_�J0dT��Ȥ���䴐"�r8^9<�*��Dh�K���Q��H*�N����P�@Ƞf���5��t�"qT�t��(�� ����c&�/�x�R����cQn_��!}SA�=�Q'�H���Fb�J�.�h���u��s:Ls4D.g e�&����WD����������	�]�r���[��땫Wt�q�Ma˒��U�s�Ç�T��K#S(��L�&�/Z'�O,ن�,�$2{����ɧ��}Ǐ�"�̀������ؿ��O}�_���-*��t��g�a��^��UA��R	3��Uj��#R"/l-o�du�P��@E747f�Β��n�)���L�} ב�cB�|�|� &����Ҋ�aY�ӯA�{8�\�3J�(s^I�M�bh��1�fҬ�����duA���p	�7][Ʉ1��D�'�G��������)N�3�9���,H� ���X�K	��JnIQ�D�`$<K�dCS�	��9�իET��B�=FK<$D���>��6+�;��A������x�����cPG�+`��Z�Q~��uZ�  �tvw6��Zhv��2�[�ϛ;�;˶�گ���/�r���E�kMc�D2&o~_K�,��=��S�� �E�@��؅�PT��ؤ�)��DV�^��o�]�+���¸b�2-�ӓS��9v���	d,	��QYQU�N��&Ͱ<%��[�j��\Ź��*T"���	n��7Ν�z�X�.R�΍��	��90fd��IsK���v���	Ɽ����Q*�xe��HH>�wMe��ղI�%!���*���٤���X��9W����\�9B�������?GD�>�߉�e~&sieW��B��53�>q��g>����G�D�9�Q�B�Br�[����8���)T8rH)*7� ��ܳ�
�J1%.��qqTT�;��x�q�u�˨�O��-=�z̏r��Ǹa
5tx����8h��m�$��v2��!U?s��D�o���񆝷.�I�ЅA�������N���i�)������L+������oy�T���i@�66�Gp����bZ1��2����uÒ�9�c�=u�ؾc�H�-��v��Ckk3^}�5|�s���Cǌ��� |
T�WS ��������3q��*�.2���}��1i���h��xJ�}�0Ʀ�u/�3)xI�����ݍ6l�����M�P���@��D[/����*�'9YP�,p&���:U��89:��L��s�PP�(�ݕNz��K����[p�[n�?�	�&����*�<�v;j#��F?�F�mX���g_ľ�'0:�G�A��;؄y�7��g9��(2��LU�!�$�]�~$����G���!����*��������pǞc����!�=�,��k�qr>�CWwW�ju��R+K ��FB2��l���M���q�Ʋ�|[$I��`2�d$�rl�s�UՕs���z��W�Q���ß�������{��s�1��Զ����D��B�<^(>���,��m��C��0���y�
�eB��G���Q�>e�d��������'i�ߊD,�ť9�03%���"���ො���@����3�������@C�B������B��?�JjQq#碟_\��-�=��LQ��3lP�4B&�hbS=�)�hrt�����?��Ʉ�:G����Vh��ʱeC�΢��KK���רS97nZ���{��r���󱴘Q�'�i�韾�}��ꊰ�k�*��	(�a5�Ȥ�b0�&�\E�~�ʋYѯ�<FE��"C���k.�Mww;�{:з��w_�ױq�fX������G��bVV��j2/��Q�Lb���s��ڴ�m�n��z�6�i�֭]-���ŉt�i�$h9����sYO�c-D�R��ann3��q�'�!�kʬ&²E����gP��?ySP4�hzzQ�ŸN%uuu��;o�{���v�`jd'N���Ƒ#�p��y/p·��)=sNT���-׷�k1�=�P�#ga�J'Pif��g�}8	D�G���2K|�N�� J3p���B�
����;U�Px�}�կ�w���#�Y�7��M�}��a�?�X4�1U>9�� ��T�"�]����p����61**Ln��,�X�FEo�մ�B���L)^�ZP���m>[b,B����~^�<֮��0���(��0V�vbr|�s�ް�FWZV������-��r���09z��!��K66)7����4:�.��r�O�H�B��g����)��=a��>���w��~�rv��Y$�,[�Ԩ$������_��D>�O=�����O�5�Tв��e1��횅%Z6P�����^�@!e�e���M��y��,VȪ�R)��0��g���[��������sL-�P�E�w ݵ	��5ҧ�}�GjT��pcS �4|$�G�b<��ĈF�ɠ���Y%jG�5�̏���"\�#�\6 ?Jb�7�뗶)�L�9d�2�y�&¦&�1=1���w K��_����Ȕ}�E��X��� ���u��#	`U[}�A$�%d
xr�s�к5�����׻�c/9P����^��3�DZv��(�����#�PR7s!�G�~7�͘��܈]4�hI��a�jQ�33s��A�ƞr�33h	G��ކDK�BV�����E��K��/�������O�")� GOLe��l��[�Ĉ�*w�?������c�� �KdN�1&�N��e��r�\X\����Pp��s��"��G�����,�	b�W��!0�gR�|�������0���;+�8���a)'��#��9r�<:{:u���.H�D7�����|�v^���_�]\�)_����49NL�F0Y�9j�y�q����]e���M�"���M3(��n1z�=��*�b^�����ۥ�Ν�u�nݺM��C���P�8�JF�+y�8f���ׯ^��;w���r{��;:069���	��c&doWON���
�����}��@KV���gϟ�-)���?����~����6�N[�ю��?iL��<TLLJ֑,ץb�)z�RAK�Fg=��-o��� O������֟������( �#� =J��45�[�����B����u!PIZ����c����W+�j�)"p'���o��^ׁ�v)+i~/������,��������,�Gq�N�Nt �H�&��Ö-P�C-��̽hfK6\�JQш���P5�^�g�Y����is9I���m�*�mI�@baÖ6�H�vd_+E����0�
��zĔML#	�wU'.b�*\ۜ���������/7M�K����(Μ>�k���@�U����9X* �]�6ױ�dӨ��s}�M���5 K���S0;������Jk�Ĭ���0�B`z�5{d�~��}������c�>��S��[*�
GQ�t�R��|TX����'Ę�p�RQ[�\��!зj�������9�8=�ϕ�hЄ��K�nŞ�W�T�apt�%�,�Q��5څ���h�\�"�@�ː
��X����dĀ_�+ 37�����X��'S^Tzr��á����ip+�籦��Z	����q�|��Q���ε�
Μ9��I$�mX�ay� N]�B��/ю�WބD�z�	Ԙ}F�)F����zZ|��JX\������ԴX�x�:�ku�}������.}	߸���ޡ[;p��pێ����NU2s�f�OJ��9y���(-��F�zq�+�Gk:�^ڷ��}���Q�192���V�p�5��e����O<s<�Sd��j�T�!���c2��o?�y\����0Y+J���V.V�/��z�FFl��O1nN�&C�4��dR��	T:�ڗwnVi*�|��o�âj"XU$A3��A)MN�x��ŲŚ˸����a�#ʇ���麀�q�UM�Ts����~TR!?FG���ъ)���U��BAl؈�}�^l�d�6?�Q��*,-�p��a|�k�P�n-(nVfI.r��s4o4n#r�B�4�.n
��������_���U�y�
�	�6�l@__�B)���п~�^�'>~��Ʀf���R����6U^s'&��bbI���4>��@���GR-��A�*�T}1�L�0����֋w8��/?�zX�	��u793)*���0~��4���ŋ�����3���l���t�hMn���)��ȏ�|*���~��˿�K$S-��pwq>�c<��Ø��4�I(��t�_��g���ؿ]�d솪[���n�QUw�QV��Dχ���OU��v���w��:����##i���"Đ�����U�����ߏ��>L��"��PR���F��XP��LFe�pR�ھ/T�ߙ��Z?ԙy����n��>�
�-���kH��[��Mu2�ea��"ی�1&h]��%]����� V�uc��9���
��E8���w�o��۵.��*�� N?���ú>?��5zkP��
7������eJ�i��7��T�Zq��{���E���^Ƞ839��h�,�Y[����k��)d��Kdd��So�ӟ>���?��Cz/ш�AsԘk>_�J(΃��RfK�m6���)�TJ�k�s�b��lު`�3�ωQe�v�qe���ո!��~�:�޽��O~'�2X��Q��Ot��o3Rm}�b��Ɣ��qh��}�ҩ��K�Š�/MOcq����+�
��,e6d�_��b��A��9����Zi	a�� ռD�,�x}9%�u� vlۂ�)uoÙ�i��Jwb���X;pJ�Ju&�[�'G��h���Gg��D���	<��Y�,,�YO��c�ֶ��?�/�޽a�Bs��b��~k��-��'Pi�9_��#MFka�ТF��U���K��+%Ůs�U�es^����'%�o�'8x�4|����x��׿�lھ�$���!|��?P��˸�=�~� b� 6n\�^���[�L����K�Z���҉�V̬�xX0shzvJ�K�%��Ä�(ѫ!B�w�hݝ]h�s_@4fSs󋪌��N����a�P=�+~��UV�<���	l�����eDs�0��s,�G��r�� ��5���0R-I��ϙ�'��>l߾w���ؾ��@�=�54�����}��� �1�)��c��=}��4�����2Mԭ;�݆��W1����@K3ˢ�Nb�k0��P��¸d�&���ӆ��7(2*���{�������T��a'�C�l`fr*j~ �mݸ馛�eӀ�18����;�Y���s�6y�PC`��"�Z�;x]	xݵ��O��;3;o~-����|JN�9���~G����� �}��1Mg9Q�<O���=��jMa�	i��H/��i���
�$K�4Hcc�y&O%��XB:�ex�굻�N'��\AP�X��8KZ��Ө\�Y��d����c�]�h^o��u� @��ɀrT���L3hx�,,�7�p�zxxP�@P�8
�Nו�-�,��U����� (����dq��x�[�AƏ�I~=ż�J�=-�1|��)�4�eG�
'�i4h���`��m*P����q����0ܴi�˯�g����	-�����#�����Ș�=�!�U�-q�7�Ă���p��h_�٤����Z#7?�<ܽl^�Ϲ�/�\�,��`��9?S[a-ӎP����kNRNOYB=�㸞)� �I?H�B�0�;�jN���ޮ���6G�''���މ��~1s*dT��v"��FŢ-7�_/�o������&e=O��@�m�� ��h *4C��,<#l���{x��0����i���qnbJ	|�N�N���� �i������Y��=���q��,��2��4%d{5.ζR"����j39%[�0�X�H��G����Q��Qn�	�y��a�j�䠆D����Q<��3X� S����խ�~�O��KT��o��'��H��عP��
'LT�j��qx�e�I�B���ylX��^�r��m������w��|E;��Ǜ��z* eq�N��W���(����s�n�p�����(�W�����,�kr&$*�>٪ɼn:<�Ƞ�M�Z�(U��l>��'�"n����J<ai���4h����(��m̬�%��\;E��͇��J�,�Y�*�*��	H��𒭅Œ�ռ�JG"���*V��]Tȓ�ɒ∫߇]����p��LYe���>�/~�:�$��¨4WLND�J�F�ϝ���<�R7��hW�6oh/ƨH�Q�6=�I��aw�ځ�����^{��+c0��c��O��}���,OV�:�DF���"�l�X$�믹w��&�3Y;y�ڂłg��8"�;��,u�F�(�^7�H� W�l�)�d%��%ݨb����8?tN� ���������$�fgMIV-�M���WI���!b��g���o��Qq#7ʃ��C�z�����e�
N���Añ�v�X�����8^� ?[2��b�A�Z���\,]O�ZF�ur�%� ҍh����	3�E�:�����9���Y5y�����6�-z6#��jl�ד���^���Jۦ>���i��S�=�4Fƨ�ET�� ���q�Ϯ'�3�6nϙ�Q����=gVN�q�ާ��,Kx�@��M���e�utȖ`fb�X�Wuch��r���7���z{�-�S6�N{�kx��I�i�%���I�!`@��M��i�����s��!__��c���`վ��KqOq����`�upq!�����2���i�c$��QD�>��L��hO�'f��f~g=� ⩴�c��x�ڨS��!���l� �O�&�Ԑ==w��ڿ�x\#��Yj~M��twb��W�3c�8?>�\9_��d�7�@��S�Zu��	4|d�똀�{��*j���h��X���9H��=��D�\F�o<Kcᆄ���q�?u K�c�+(/��r�>�90�6f*��c67�{ٺJv�Eǚ-X�a;��$�$��j>2vR8�Вy@��d���a<��d�����v�n����?��Kͨ|���?w��9$vj4��h�>F����UL��V���n�U�Y����Kэ    IDAT�i��M���N�8�뮽
���8t��_��O%12>��[������@�-�J]#\l봦[����g>�y��IU�I�,W*�y{�<H����6��̒�f� I�_,�p��)�ˇd8��TJ�0�G :�8��޾����"�j=�`@�Dn�RퟪU&8jò6���8�f=)x�E�kQA�F/�"����2FG.h�Z-�o�U��i��u�]��e7�̔jr�����Ο����[U�.&�35?�K��y�1'�5 ��t)�xHI���a���z����+���l���f	O��,G=w����F�\u��"�=Q�+��;��'�..���kdk�U,7=�������G�c� oߺo��_�=!MN ���p鎝���[u �]����խ����1?45�`:��MS�:FG/ ���;c߾�d,����e^y��tj��Bf~Q)��ba���.$b��'��;���56k 1���U8�	���o���34-}�Z���]s_9���yc��^؀�����<-_�{ӧ����D�r��Ɠ݁��S�������G���x�8�.�' gK�b��h�E�,((�-�*��
���=�Ȫk;H��ܲ�#La�AZ�ӱ�&]X�r-�YJ�[�aȧ&�=R�5��^�S�T ��sE�|𽗥Ii��g� ��6^�,�J`�x�X���
����Q���؈�h�^*!�R�\�x\z���I�A���.�-�D� �eH-�0K=�%HeZ23r|��P�C0��x8WWw��3��G���x�j/����
pi"�i���sj8xm��'�w�YI��;���9u}j	��M����sl\���ߞ)�[�ϸ�u��.d�x�Ο���|l�i����Sj͸��׮�B�ar
Ó�X*�v"��E熝�:$���,|�H
�O�
ũ$k�}.�(R�����{XXX���a J@���>���W�*��ժ�W䣒_����y�N]@��u�~v��"��y;E"(�@�Ɏ^�t�AK��Z���Q�Q��I	�����oM��ߝB{�/��g���}��,�
 �(�n[������_���?����g>�o�w�<��g�Y�(ǌ+ZE�H����߀
����.g�ߛ�_�*�3}�a�r˫0=5��~�{2^���eT3�0�^~3��9�/}��*\,Bpф�`V-_��4�ɼ�ЈEY�����Ӛ���~�E�e�ª���T� ��Q+�P�%¤�1t��!�,�Z⢣����r�i�cc +`V"���a�M��K`Har��(XR�'=X�I�L�TGU�kE�N�t���0|�����ɍ5�qj?�n����p�׉= ;��E=L&���Sg�O}F׌�'������PY�Op̊;H�p�y&�֡�t��W@�T;F��rv[�����aR�����mX��_#�;wmצ�v�:����q|�+_�YR��"�q'����^����
�����_{��w`��:/ A�@W������^��Wir�ש��� 9��
6���@0�67~���,��C��� �<��#_?�fyHP�ϟ��1ˆ�\�f\��蹶R����YXDA,���n��,��+���(g�{����w
��Gŀ��ekq/�������R��?�s�]cO��J��q���'�R�F��/T���P�C�^�&�LD��dG���oE�`� �*yh��!�KK���w�M�z&�k�3�^�?zg�z�Ꟈ��s�}ɖ61�: N�&�NXV��U*�����Z~@�SZ>?Rm����u���<���E	�����"�/k��-�iFr��F�����,���n,Ӕ�� .���]�v	�]�k!P����(FK�9�h�{��_>�z�^�yOh~n���b�~�����w<�lY����~��Y[��L.#�X����Ve�>%��uD#�aNۇ� �� uPf���K��������F1|~T-�`",gZ�����,�"ز	�_~9������L�Z�X�Uh]�N�x��>0�a������69�C0@p��Ѧu�B���@E��x��!�3��C$�@4\E�����gF1?6�J1��f���r�& m���޳�k�!�n��4�*j�Bf��$1�F�H�XݙD[�4r�0|{�Bn��_@e����>r�o~�%*�:8s���8�]���)��ix]�Q�Mz�L)i���}U@�K�m��7ܪ�[��\u�5�b���у�`��MB�<� ���nǅ�	|�_���Y�g����;Ի�����s�Tk�Lpߥ)��IcT|�&��-H����T��m��B��H��2�����D�
Xɪ�!o����%d��<����q�s�Q`Nl�aq��M�?��Sp|�N�D�T�S��%��iK#����S����{��|<��VŚ5�q�}����߈�<h�V��d�cGOH��qU�;������Z��X+�_z�7�_�����_��2�.]Rܦ��M�/���R�6��=����C����F�VA�������� N^�?dQ|�p�B�^��5Ǎ�a��d��0�p��a�\��J����^�:�|���s[[����<'ڌj�韒�{Ww�6���ϪJ�r����\Py�G8~ۭ��-پ�K��M��{�i��z�|�{n)#�B9���3��hy��Z��U,K�'A����T&��v��"�5�)��ք�����B�^zbgV\{�E��%�,�]�zfa�~� ����n��F��&��1"�hme�����31.7t��p4%0l4i���B6o�
��Xgr�č�S��-:�#���$?�P�E�bδ�:PI�Y�h]*�!�J	DK��	�	T�2B�:Z�*h���Z��D#��o ����!˺R��L?��=�o	T��ɢ��Z�����ب�PJ�MB���!<��b������b�rq�a�þ��b��w1P�mHк�^�W<���s�X'&��%=|ho#6�` ��l�sB�T���P3t5�7���R�M��3y�}#�I Z(D= 0��v]�S��c�Y��싡�@ у��툦���
�����hWN���F�o*bTTf���aAB��盀˓�e��{��6a"@"��O9�_!��A��\w$�<����u���$@�!_��t �p�P�'� ��x8�X$(]Lw{�1��"�O�����)���#P/�n_�v������ڽ������W<ul�#�z��|���+�0��q��̕���ԫ����7�U��L�p�^�F��/|������o������;���}k���e�|%�'��|�|V��9d8��oP��7�&�U���� ���&Pa��W���D@.�
iq
!��Z����BnPdS��T8��ֶ���%☝����$�L�%��C�l���&7g:jRƳm& M��M1���3��<����X����$#��m�Z��3�ջT�H���&R���Ї>�믿V��;�s�E��_�����Fi��u�����4(�r��%5���V]�% ���~���W���C�b�B.~��BH����ګ���)+��/�T0s�zz���O��?�xtE��,k�����Q�fD��/ �������A8¤�y��nz�%�4��fȲ�V8���(n�wrs 0�koooՆ���?ŷ��m��r]��`{Q���١J�t���J0la�j�0'�/B�S<�͇�Y�Ĭ,s��r�^�t<#/�i,-�v��߀TK+&'f,�� Ntx���y\��i�� �dh��m�׃�����N/R��,��AT	T��"�&��1o7-#�Q�V�*�c��d��2|0}!�S�J�W=��~עg!���o *t~M��/w�Ȩ(���Q!Pa(����i]h�ȶ�*l�0��_+a��^�Ȉ�TR���)�����<�C���bp�"�@��[�\C�HL@�T�H��@PWFV��uF��	� m*3�����P��s��2��X]b��i���uk�W��5���@�.�"�Nx�y��9�Cj�2*S����c�H�#��c =�O��kQ�!3��h*�L!�:3���-6
�,f2�B��CŗD��]h]5 FEm(3ˌQ�d��\ٶc�� ��*��ZP)�]�G���A
�)w�u�|��[K�c�Y�r�9�Ӛ��;�!�1�1v?�����)��ˬKa���*�Rʰ�Z��SC�Vs:FOG-�:��,Μ=�}����%�U��ȶ�����w����o�~�G��)���+ֻ[���S���Ce`pd�"A*�)���ەƫo�Q����s�bj�\}����+_���X.�l7��j����D���[�Ⱥ<���tww�����g@U���&M�@�<�J� ����=�f���UE� V���7����ǳZ[m���͠
{�S3�%��Lq��N�^���(�l�;��W��󛞀�D���
6_:	rD9Ш P/I�B}J:B��P���~ �b�������M7� �-�˘�YP��w�G�3݁7R����G,S�`�UXN̃�Q��Z��"�= ��
Ϳ"�m*�����2͵3�ZeU�����v���2���$�l������W���������A@�ﳀ��,;Di�E�(LF�BCs�U�Z< ���2���ݣ8Ntw���a��hdFlkAL7[j]�'k~^�:�i����6Q�\O�ta:��E1|v8ޚH�X�!���j�g�2<��XmN%@�q�/^KC� �$|�Al����Ĵ���$�ςjCu@Ž����r@�m�F�����_~���F�Al���ki*�[����k��!+�� ������R���=��_�$[?*<ت���	 ��+z�hpw�:���ĵ~~.�B�T�AF�b�BFRץT�*,����*<Du�e9��"!?��ucUw&G�0��`$����C�����"X�A�	�en�LK?��- [(��`��WIS��/��Q_�vf�~�m]�-��Z�+��;,��k�.?��roV�4��^8�|!�1i��[fzy��<�}�9��!�bm٘Fu&�Q,�R�l��lu5�'�niA{g������X8��|"�"��a?��Fq�ܐ������6� ����X*QPۍD�z���ˌ��L�Z?,��F�Ľ��QU�\1����1��$�Q�+y�����3�������2�R&����>��:c�g��c��W癠3æ�R�:��AZ�hDSg�"��ޚ��V$�u�K8q�0=�� Y�zadǺ�O������7�{�}TM����|��K�*���(�RѦF�B�ʣv�>%L��&X-�^�a�v\wՕ����(�ⶎNl�2���ǟ�ͼ��+p���cxx����Q)V4"V��Y�ԯ��[��Ӎ����cpx���JC�?Ć���-���yx�n���aEC�_B�C�� {�i�Zv����6�`��zy�5e����9K-dU�JA@�{��@0"S!��� ���{��j3rLU��L��A҉|��2P�ţ���@��5�Ч�յ���k�uzz�N����.,Ba�i��⇫�y?̻�����r�[7�#-��!��+V�z�G�F%��m\ ��q-LQL��8�����C=�����߿Ǐ��3{���83�x=0�r��0ѩ��q��N�_�L$<n
8)/ID�����3��y(��H+j���a�?�,d55D���,m�3N%@��S�����o�N�i|�U"�5�FMp}�9���Z�V������N�#?��� ��Y��1aU�d�֯ۢ��щI�J=���nrLn>�{��Zb^F��;����p�օc�� �4B+ڊhWk�m�Wk2a��&ױ	P���v�j����3R��uu$��jMkҧѐnIc�ݯQc7����eF_p}7�~���*m-)1*�F�z��P!��h��(�U\�y/E���/��*�U;t��bQtu�c|tS�c��QCEӎ\�d�8�
0$�X�1>2j�6�LӅ{pxX�8�EB���@_����d������@�P���qn��Z{������� ��D��e��|di�853-m�_��3��rI�(�j�Om�|}~�tuw#�jS��[�X��zЗ�>Y�H ��S8?t�Ra���jr��懭�s��J�B��?ޅX�:�m�zdR7������q�2dҞ��hmI!�0���)0�=�caz��C�FQ�GS���ƈSm�x\�Y���g`���r8��T�l9Ȭ�4S磽0đpk��2���tE���T:�ގDCu��ǉc�p��T}�6���;>����_?��}��܍?}�Ƚy_lw�},��4�hJl���U�yU�a��H��$"D&��p�U:��-�ͺK�V��ߏm�v൯}5N?�����*e����B�P��q;�z��}٪� �uC���*K�(^�''�E�gsK:�x�4�n�:�d`א6�s�T���S�x��
�G*�\�;�b�&�sG�d,Ν48�؂a�<�l��wfa�s�d�(zz�n'�e��&���#MKBk�гA�S�����(�ڵk���N������d5�Ǉ�l�Ԕ���`�4�;h�i^�Ǩ8OV�-ğ�Z=���Л����/*�4��t>�+�(&�҄-D��2>�7�φU���z�w�RP��[�tyu�o��@D}}�V��IaE*�^���M �����и
�!��LZ2�`J�qdKy���1�Sf�l�n%�5�a$Z[$�T�M���P��J<������)��```�����TS�9�E�D����q�&mD���&�.�t-m^N��Q���x��Ҽx&]��͌
[�5$��3�+nV�JseMGi�Jr?��l��0�5��ƍ7^��������=��������D����R�Y��1@o"[��?�@|�e.GF*��J��C{�	T�R�.�R��@fi+�@�֑ho���zb���	ںy^��15v�������~���/an~Z6
��b�r�n��կ�W\���ޅ!>7,�B���K�\cʃ��h�����{�9I耧��aO�����&q��hֳah��?Ǿ�fr(��������2hc�1�s:������@ YPj�e]�{�U��Ꭺ�6[Db��1������ϊG�����UX�̕���B�0h"A���DRj�o޸;Tqfh��"ֶ?��k�������
�u�x�𦏓aE -d�禑��F<蓮sl�.�9
��4�4*2��P�^c��IV��p��-F�����Y"�4��o�?9E+0�	T^CB���,��pO���2A{kB��z�����c�d}��h�Gw�k�����x�-������:po%��2_����@nQBj���KDh�e�o�N)�S̋\������|�Z_��W�����?���	��Iҷ��n�������G�RW�JGKZ0�UW_���^<��#8?2�ѱ	�WVQ���)D�A��5�%%'��b�˶O�f`EA�
��6}cU����Z��/�O�z���X�ժ���&������w��+�J}��F����I�=��^K�a�J5ԧ��v�P�]Ρ%Bc��9�i	T$���|�ҝ97I>�\�	NU3=���-mJ�&��C�n�*�='G�J^Ez�e���XE�6{1k���8Q��R��TM5oX�p��1f�י���s�OK[OXU�M��<:�懴>A�=+*�FǨ���n��C-#��p��k�Q_čK@EznbPXf�TDT��S��RvɫN2u#�̔m��r pI��W�HT	�!f�ߊ<HM\�5���zz����ږ��ٳ���lkU\)�Q� �咜�G��߄����i�6	�g��S���'��#�cA���$�{�l�}fx��%�ywy�}�D�M�^��u�F߱n�j�x�S_�k�{�)g*�<l2HOk�avvZ�vw���N���}�    IDATJPΑ� �*�W
ּ�\�Q��։���gD����BfM��M�ʿ�hl���hY�-����yFx��(�{��;𪛮��S�q��a�MO�@cd��R9���9E0����_�շ�Ζk!�W�؅�8}����cG����/.axdDU=�HT��VŴgb�<�S��E@����p��{���+`���eTV��}-�t�t!޼y�Z�W_�G�0�P�I���'�}H)�f�g�sj��+�Xa��*�B�,��N$�&ŀ&R6Jv��gnzF����e��J8QVǂ�����Thmqrh�x�k1��#��A�s=B�T�*�92��%?{��ς�@��fu�՗��A2@�W���Ø8y�d� uh�1�৾�Š����nΑb^g�_�q*]b�Ŵz��p�A�5�7^A���)�e1��kW���O���5.�d�D>��N��G�F~lWǧ��=���k����h)�ܿ��9�~���5�d�=%�J��kY}V��Ҧ8GAr"�z�C��SK���[:Þ+.��>�7�I�?VKT��`�������x����5����[/���Mp��R* ��J���Sg�`%��5�@3&_͏m�XZ��En����/�R� �z��"�P�!P���5Ŵk�V˲������0>6
���T�JAM�syq��-�;{W!����m]�������.��/؜��N%h`Ug+*�%�А��&@[ty�x=�Zb��B'F�u�`r�oU/�����h�˲'��z��@�&�hEU�o
�p�YP��k�=ǰ\J܆�~�ŀE�ff��k�o�M|PD]�����9�X(1̒c��k[�e�R����j���INHx��*.������V�^ҭ=�&6�h�Ǽ�|8j\L�5x�0�=���VJ�#e��E[��דU-��w��z�<g�s�Zj�`��}96m^��<��4)iVN!?ggВ�<���C���������vl��F�L`~��Y�����ڰ�P*�Į	4��7	���uV������YSk��Ck��Bc�MFpN��tX��ɝk-�4��VH��e�+;������G�������w�T(��{���>�1d�9��gs�AP��T����!��Z�Y�Io�ĜK�~��D,x��WI��T���PLK��~��~�\+İ�P�^0`�z��_�	�iM�3�Z�W�ځ[^v=O����Gq��q�����ӉB.Cv�<}B���5�d|��׿w�y��%��139���	���;p� f�06a����Y��z-<w?U�{z7�Fǎ�u�tv��,���EN��p���{3�b� >1*���i�=�W���]��d���3Y*��Ƭx�E��\�l�P�AGb��P�����zq/��Z)�`<_؏
)o�,���y�FlܼsK��?މh��9?��Hum�?�T1��n�ƤX��<cju�丿�:?=�Jv�Mz�;q ��g �����Q`E�(��3�g�؎��g �Z�����ud�jX��Ec�1�*�D��M���mٲ	����H����:�<��=+f8�QZߵ��3��߹o�־�������?z���j����U9 �r�"-K(K(@�hT�2}t�qJaIS@��okmA�X�А��<�H��a�\9�-��U������Ƅ	n8�ֿz����t*�js�'�jb9�&al!��$�Gw>�m���P��d|t�sS�`���Y��J0���
2Ej�x6��&7���޽{Q+S�P�~ �E]�b˖�x��n�ͮR�Q�#�����)�3�#�Ү)�o�?���8|�Bո9R@�騰�n�J)�������Ν=#FE�	�'2���	ޛ��hנ��*�4���*i��X]���m,N��6-&ƨ8����d�	;R�
p�/^�͇�l�=�"��$���f��؃�	�e�N��+*-��<��*�>zE�(^��Qu�TXӪ8����@�Q��)�"��m\���10f�,\0d�ڐ��S����U-mmF������ڞx�I�%�|�=Q��`������7߄�{T����$ba�5����hoiŎKw�w���~dmj��K9?~>�c���ٹ��׹�%d��7a�矱l��1W�Th@ݻ.+���U� ��þ�g��|x�Hhc�}�p@��$n�L����ވ?��?�z#P��'?��lݽ�����
7p����*���[(�!gk�%�X�=�{�"�zzP�FE#A�M����
�V������H�Qi4$ꏇ#س{'^v��8qx?Μ<��1��SH�⨖���n�S�<��@���n�%�q�:�������CG���߻��b#�J�'��7�䀧����2�V�xƞ�������8�cK����;�~PqbZ2*�."P!�A�If���h�P{'FH~@��L_,o�޻�,��ŵ�(� �dK��{\O����?E��k��4�d.����siaC��*�t/2�����ڽ�0Ź�� ļS\Kwp�-�v0�V�T�*3S����4@1~��&/ ��9�a�R��S)�Ո�������J ��1_B aA�
8TA���n��+�5D�%����2�]r�%ظe@:N�ѡ�����{q��9+�8%VΎ_����G��e[VYv�/��cT~xd�����B�}��j��f$FS��x���i��I<,)
�B?���b>���sl�pa�ն���i��4I���Y�"�B�5�f��G��	X�@�ZB��S_��,�IgҾ�a`-���F(H��Q�<D�� �[���'17;IDa4i�oZ�{:[��>��ڵk�}� y�!ģa,-̣����\��JlڸW]u��S[[��~�V�泧���{�ܾCx����$��۰	W�p�9<������d�O"�R��!	��5�r!���A]3M_���縝�0�A���@Y�z��q�h�o���J������1����V�'�t��O�!���7��{�I��f�}�/�ު7�Lj�-���q�I����t�jt�^��ɲ4��M�N�t������P�C��U��{��V���b!,��F�<'5��B	�=�F`ž�����H��Sk��]8x� �<�MB('���db����I�v�/����ajrL���x��y�d��:���\s�5��?|���fKK����ѣ���ÏadlR:�|�����KܩgЁ��m��8��o���iK�ͺ�XWy�k�t���=V�{�|:�Ȩ���P������wT��׮߀���)�6LdYU::�C��:��u�9�I!P�g��/3*�C����iڭ1*�A�@�"z^bf)�׽ZSGp�έx�[O=�S<���FOG;�{:����lų�=��om.ٶ��[�*���H�qL���ؑ�z�=�_���l�#T��0�9 ��`w�R��g,����Ĝ����S(��>�V��ѕ�I�s��0�:'d�F��*W]u�2������ �xn����G?��ir\V�]nz*90zC	���
�x���~^Gw���/�b1U��"�s��(7a����
5*[�l�����4mG э|%�t�F��^Td�FXb�N��T��qH@����Ks��h�F}ڒi}5T�I�������G���Π�!��E�A��A`�x�(�L�Y�;0�(�[�Cv7G(��~�C0��Kw`�����H%#HDy0/�ٽO��А��ō����{���?~�G�x����&v>{��'g
��������2�#��| ���z��J�/(ǊY�UD�������4Wv��"�D��g����*uQ�qXy���)햣��t�+f������]Rs��b���%A2�y\>�J�#��J3ҝ��A��Ј��`�U���3�؊-�7�����8�ޞN���/��:	uy��U�B�m[/��uk17����%<��3�����ΝG{o.�s5�8�}GO!�l�F��d� �<J�9t�b*���ΟWK�2�BM>32�
�����ԯ�b��Eh�h���+A�@Ř;\/fT�Ad�ıd=<�'��p@��on$U�K �vƊ��;7��]��s`%Pq��P�#�`llD>x���#���ʞ�Un&J洙�~-�:*yM�Z�/2F�snU��by����Q�
Uo^���Mx-;�h?m�Rl��|w{�Z=�ݽc3��j4��	�P%�C��ڌ!$�1���7`�SO�Q!HFeav��ܡ�ߑC��Յ[_�*����=l�d�6��܌�
���~�i��cn>�\����9��S{�M��y���c�ʱr1Pq�Wu������،�\��^�Z�a��wN�X�O�[B������j������'>�4]�0w]��(85!�*�2�H�n%ixk��u1+�*�٠K5�+���`P+�@�/*<���]T~x`𾴴�jϓ���b�%1!k�����-�bzr
s3hM%��Վ��qT�1:*ժս��������Mo��I#ƕ*F��q��1��ƱcǑ/T�8��͡�4��̳���wBq�n5'i[��ĘU��'�/'������*��[~��M���#�~��W�QaQH�
���������s�|\òx��,�ɉ��ғ�bS����������@�%�)0%��J��C�-�\���&�6��Ǧ-�qa|
g9�n�("�����X����~l� �� �*��Jf�rN�"TlxM�<�\j���m�l��z�cQ��@Տ\6��K?>Q�nb�D=�L�<IBAf�d��g�s,N��ظi=:���K���K�y��G1<:.=�������]�W���ܰ�w���؟���'�/]rjl���+�� �T���(��8��Ƨ4�"#��	�T�)� 
�E�\��$��	`�e�����CI�5��cS���:J���z2���Ţ�!dUH_��p6돳�&��>{��L^=P͕s)��r1���)!V.��r��K�zY�*�+���nh>��kVcc�Z�9uR-�t*���kny%V�t�aP)�Ap�cf��7"�҆���c��o~ÓS��?�*}�9�8?�&�j�196�@%�A��P�X>3/F���| �pJd�m�*�:��lWD�Ν�bpp�A2يΎ.)��x\Kˉi��1/6��{ǽ�ć�̸,��63o��#�u�~�ſ�'���S���#���a���-����%����d�s�V7�J�r��W�j�l�]�g�C�ME痍3R[��w�Jt�k�_��U>#�d���m�+9�]*Դ�I_s!Hӵ�&�X�[�rX��N6
���rǝo�3O<�3�N��K�#�.-b��2�;~�:���7����wb����9,��cpp�<�N�8��\����j�:�jrR.`�t3Pin�9��43*�\�Q�ߝݴP6]��w��{�H�����ƨ�Pa!t�u�����Z�� ��G>��	��s�ƦtXɳ&H_�0�`��NR�:����� �0�4EئQQ+�V�v�*����^?2*����*���S̥ěrp�v��H�'��d�BcÈ�CX�~�G.`aqV�&�޾�G������^�f1<4�C�X�>�ĉ�(�jP�9��H{����V� J� 
��aӡx�H����f3Z+U�3��z������g�����>ŏ��;���S\��*|f�론~��
\}��缘���s���&6����&m(�&���]�kEm���lN��h!���!�T� H��P��q�F����4j!�N��m��@k��#I���~D�.8�2d�g�\���B$j�����K�*N5u���4��C�X�K�W����Y��v~Ӽ��J��W�#5}F
���}��������rN��KE"H'izC�_D���ǟx��3���䫖�ع�������G_r�r`�8�P	|�����gk(�jX\*�%�%��s���>����쌴'�`��yq�y��l��U����^gۆ:��+ET� �"�)����^���I�7e�V@�"�A]/>����3�RT��O�Nhܫ^D���֠K��~]0��2s�e�g��X�7�H�c�Ϟ:)[V>�T����u�d0?3��6���Q"3Ai�m�w!W��ѧ��;������oy�����*lP렱���**�%}e�����n�2>:��V��6��"�2��z��W�B��--)K����OZ��?(�7��}�f���9�6UE�m�&
X�hވj����'4t��J���Fo+Z�114�JQ�y~�bSZ�
��r��mrw��CL�,,��T�E�:hr��2��-2Ӳ�F����BE��X1Фl���tS��Aӭ��3�/+C
��>Lk�ƨx�B���hk��&���&����ↆΛ�+�b�HD?�����{�܍�gN#�YкM'�j����j	����s���w���X�q�6j�����T~�;vB7����*(�dє0��Zk�c�v9`�|�4kt�y��$�o(ˣ�~�&�������}�A��ӥys��3C)�}�)Q�������򗿌��ʱY�q �٢��Ξ��l�a��m���<ļ5�C�c�dɲH��޽�P��
�<�'Pin��Q����ե��z�7�P+��5����.?$��R��qC�����1��^.�����[���'^�R	�����j�5�1*FF�e��髬���!y��p��x<��S{�����90C@جk����s�����"�馛4���&l]]���Py���u�9�Ip��N� h�9��HD<�ҘsG�*���sR,b~Kd9����H!����"&&�Q��]Q���v�ƍ8=tC�3(�H�<T:VoE�}�2P�n�"����Œ�N�9e[gvfR�=r{���	R��M�t2ͣ�]D,��Z*yM�0�S<��$ �'R�q�8�D�\��b�r]6�P� u��HIE"QH"s�( ���G[K��)<��#�Z�3��� J;�u}����{���3��0�+�cT�-������#�����v.1�5��q\�F�ꓨ�6�dԹȹ�ʫ��GV���S4q��{Џ�%��dNL���dC�*[~�P&��BQ����A�X7���%8$ �K��s����FmF�XBXbM�6Ҩ�@�q�VͲ�/���Gva��j��*e��I���۴�CgϨӳ%�_z�kv�`8��u`�
e�^���I��e7cݖ������ڋC�"v���Wb�ѓ�0�(h��*T�u�(�
֐�F�-�bns33�!be6=;/�����kV����k��k2�G�P�����=FG����}S�I�Q��X3S<ھYd����G1
�z��*�d�(���:��i*W�͇�U�VٛC����߸���Uuδ{��[������_��S<��Am���\w�DBߟe���1*V=Z�|��O��pO�-�+�)/���X���ڤ�������B51ho��Z�s�N9�j�#@�Yӳ�>�c��#�>y1/6�D�L�V�XN�Se�/A÷\�̒�3����w����;�z'�֮�*e2���TT��O=�Ckq)+�21=����Aըae0b:�E���}��׉i���*��*r�k����M�`�@��Sn�~掰='�cI��Xm�J�E���n������J\961�H<$a�=Բ)d��7�K��	�r�G���������y��������J��F5
��b�5>�i	TZ=FE�c�&M���N�j���U�57;m�]�{T��a>5�wv�0�;ށ_y�[�'j�U151���<���,F�G���Ads%�NyFRxf�Z�^k������/~.u�?<�	T�^���7�b�}�>_tX9�cT��2aY�>Dւ�
c@PY��O?�>���?yX{}Td�@M�Z7���>QkWfk~�M)�-��1.*�,�WTT�8ADc1�N�����F��� .۵����ĹA��̫�S�#�\��5[Jt @A�E�
���{ܞ���(Y�'����BfqN�U�)����ĵ�i�V�dl�QD2�C%;���v���    IDATT�Y,.L�V��Yp퇣	��w��&I
�钤�(�������2��Z�R�*��DJ�no�#�"(#77�'�|sٌ�9�Aj��w����/=P9<Yܔ�����nϗ��[v�\�ca>�s����"[����
������ng8��Ĩ?v�<[�	j��Q!<��
ָ�g�C�\2�B!�SO�:���˨&G$S?nll�3�=Ҿ[#t{ �� ��_Q~*���S%PY@v~��ꕂz��T��G��:�156���}c����M�]�C����%�ukנL�HL�����Wb�U;��<�/|�[x��}x������atjA!Q�$5�V*#�V̂��W{2��Ҽ��Y�WK��N�:2*�~����}��4=$������c���=8{�ܲoY�[�Z���＇|��cUV�(iuS3�m��/T�q���Bq3op�:����}}�dhG���[�N|��	���%�B�@���mFjȪY8!E������o@گ���v����j/�΁6�?�]�P@#�b�291�d�6o܄t��<󌮭���g��GQ%��(ّV%���FF JN�0]���cxhP�2!SoW��N��= s,��r6����p��!<��^U�d'�Q����PH��/b��w�}z��־ׁbg��H	�V9&h��o����o ���PD�Asy&��g��d������+��ޣ��مyM���h_n�4������6�@�����DS���ii��M!q���(���|M��ڐ�1ٷ��-�"���Ҟk�Ǚ�Vftl�P'U����c��U��j����@��W/�����7,��"c��8s���ف�L'�n�:��o�&����YD_���gf��޽*J�GƱw�>���gfP(W�ܭ�әQh��V�:�w�[�O�a��̪ݜ-j�D����ˋE?4=OJ;P1D]]Bfo{���u�]��O�k��;������Z3�<�� :@ſ"'.ctz��]���"��M�Z�.ᘵ����p&�f�����-)'��#�qB��F�񹬘�:i�P	�:@��7k��~f?[{��	�5��k;=3!sKb�)Z����|���A?b�:�sS(,Lbz�,2�#�k(�� _;�6�.�bdt�Jmm�����ѽ}� Ncv�����$*uQ�b�!Ƣ(�C2F[:�TF����ӏc��2�XWZ8�c}����O~�#���=�2*���j�/~��޷���v�n@ ��L�Nc~!'��#]m�j���otdL��F�Y7&	S,g�a�0���E��Td8�mԞp̒7�Fݯ)�b�l�&-�M!� ��gYbD�J���aiaSӓ�W�2m#�I"[��Ч�-�h��؋�,L� �����C�R����U]=���U�)7^{�Nm��<�y��m	*(l傼��UU}�����o~�N��ͯz;���FQ���	V�N T5��і#)�jrjB^.d��cT(���?x7��v���:`���D�3�8u����������uix��s��p�����e��mJ&�s��D�^��g�)��U��m$��.~� �F����R�c�ɻ�~�����*�ttv�������?��}R�o�b2�J��LUfD>%j����Խ~�7�V �b���B#m+O�B��N��*��$�f���{�(���JtߜS�ʩ�:�n��Ȁ����؄lcl�a�`<$L�1��6���~6&$Pj�s�NUՕsݜ󛽿s�J����1K��V��+�{�w�o��o����hԪ6m>nB7<�Z���~�;���xy��B6�Z���C�-�'�X��kB��n��2���Ud�)10{�A��?����}عw�b�91q��gΞW���naI�lm��t��ֈ�8%���>m1-�3n������Y��ʅ��o��?��B��Ϭڐ���>��7�[�\��̆�b���w���u�7�7Xc��A�?&�t�<�3�{	R��S�����(�Y������ql�ɖ��,� %p�=d&��0���h��OZ�S�]�!����$�r�S�b��H`Pw�pE��j��һ�ާ��� �g���� ̀�J$"F�o�%���o�!���;s�|���2~�������ͨ��8$*�Z$d0�������Vaa���,[^We1Sǲ��������|���k"�ȑ#���������ʕ+�����=���d�G�:�2�n1 <��c1i�ĳ�(�ucrn�غ�[#��v�K���=�d�y�>��rG�v���I���Ҩ�xb�H�'��x��3Lm`��^9o)��y��3�♍�J�����u_'N������Z�,�&�"���j~C)��	t/y�At�&p��µU��@����'/��9t3z�w!�ՇJۋ�\����U,	�z=p�Zj�ăNtE=�X_Y�S�<. ǯs�_��vhwߗ?�_��;��g�y*ә��J���'�\�{BѮQt\>,����XD:]4&>7��Le�I��l���Y��6�G�	+U
f� ��{5-���j�f��N�.�&���lٗS�xnޤ�)�d�H0Ak6����5K��2��<Le���dk��ú"6��4��VL#���jq����!;:�si\��'����F��p��sב۰cxH�2�v���g�NTJe	���م[����2y�)|���T��÷���".OΣE7S˝�@����U���@4��3-�VW���5~L� r����o�&^��WI�-�(+�fGt0}5��/��S�p%|�������M�I�]Im͉�Z�-�nj���h��,x�_�dl ��J���ь4������N�w����r�e���߃��$��p��$>���w���gE�e>9~2ȋ�9�	�*�%��Xc�J��gĶ^��7KV��su=e6f��1Él!����ܵb���Y�Cv�/��������������*
C��R��	�P��4UR@�� �E�,��Z�PM��{q��a�sf�LMLjڍ�������:��r��˞�2��- #�j���#D�^+��2x㺡���֨J�V�[�Y[>5��~�h3l�FP����7{2�>���>F%���dr2`�m��D$����km�?)o�,�׾�WfД�� Y#�6@�V�fT��<>?b�J��P鲀�a�l�B�7>M%P�ǢrO.3�*��|������i�\Z���g�O^C&��#-E8,S�_��_��:G!���)�q<� "�ʈ-�V����Q�o�i�8�)(�4_�|�V��LD��2�aS�$��2ƞ�x՞��	��]�l�����/�)��da�$˿��ϳg�bn~Q��/������ ��m�r�S�mY����{�60cMұ�uZ���}[�&��^�iy��#��p��4V�5ԝ1x"��%Pq�{��F�Ztz����:0&�|�b�}n�>����0�f�"�.	H�V	p���zn��,M^E3����	ڬ���MƱ{lw;�ŕ9<��S���^����gΡ�p��H�o�>t�B�E��h3�k�o����L�;��T���"�?�2�Tc��E3�����_����g�;г����ʎJ���K�+oNZ�`�-g���__A*U@���)�B��.�!l�lR��u�[K��r
d��T����77���;�8����?����6�_������/D��&���9�@fc}��0BA
4���޸�H�Ň� D��[oT�(��P)l�S+�|��%�]�#�'0s�����`@(�+���e�CovzÃÊ�fN	�O<����'�/�m�c{�aq=���4x�uښxP�e�.�B�'�yv��z�+j�)���dTT���w�g�u�s��hqd�)1-}5��ſ�ĵI��Px6�bkT؃����vQ��YU�QT~7D�+R�[�ۙ�ؠŮ��?7�]"Gsx�hZ�c�d�V맿�Őai�L=�=)�ԧ>�<���8����C'�ϙ)3	"y8�"�7+K\���~�&s�	?@q�ƿM�Gy��+����,0�����h5M���n���t�am�)���LF�5*/\Д�(�)��b������5�@w2�|6���5�h8>i�����#Q��&3��X==��ҁ�����"]]J*�����=P����rw�b��6��t� c{N �a�:3�cr�`�Za[�l��0����5$�fԅL����x�_(怾I�w���en����&P�z��H��m�"FEkC�<-���@��6��Ѯ���4Z��p��g�E�Z ���Z�j��h���c*�fS6X� ��p:g���d�T(���A<��+�p��̣����0v�ڹy?��Q�P�7�~v����	`r��m����"Z�c�)1wk��v�6i)ln*���Z�?���֏����:��ֶ;���ũ��	da��� O�9���T�O�.i�l�"��m@�%!�4��o�vm����=��s��!������*�p7B�#��wp .T�[��>�'C�ԥX��	��d����MF�,��v�m@������Q�.b��IT6��Fq�A�����>�߷�h¡ J�<
��=݈'z���.^��7��|	p������=��v �R���z�;����$��]!��u,.���Ǒ/TxDyP[߿�������|���/P�JWF�u�����K��Z�@���c-����Ul��P���ˍ�d�����ӛn���db$�Z�YE��C�R��^�f��މ�5�Ç�� ��]jW<��I�����y��r�(�M���:Z�o�-!�M[h��7{ֽ���8��(����^*�Z��2J�1**-DAt��XYZB�B-f1�^A$2o/&'�IC@-	�{VA<������3�$Ȋu����19���u��r?%P�S/Z5x��R����)
���fF�;J����~�WE9 d�9����F�y��������-ž�L��fQ��5*h**�m֦��|�sQd�����T�?+��j'X=i���7�M��ň��w#���C��w�y}���\*l���D��[�&������'�i�-c�S[�\p����J���c��l��<;���hS$P����TEG��
}aiEp]�zC��+�B92�}�|z==�����V�T�fLwfROB�kiIZ�|,y}~�z�p���������R���ӓ���/^7WۈyY�f���70����,�N� O3�Ѵ4��׶֏ͨغn�*v�m�g���e"s*/#��Ӟ�^(�5%h�o���i:���6���Alc��j�Q�N]@4�Ѥ�Fz���$�ɲ��D~��c�fnSNrY(<hY�xMQ��>�=k�P��e�qT�!�C��0�$�~8�(�m�o7�*���l��gā�T�3*͒�cY�ʘ�
]i9�s}�L*��*|���i�3�+��k��I�ӧ������?3?��A<��4m���E�ޣ�xuج���1�[?�;����.Tn+7�|�v��Κb�%V[� S؊���ͨ���$��Ӄl��׫}��ːm6��j�ڹ���v'D�zY_K-��(T �;���f��o��&P�E�öi��h;��eZ<��P�ŵ�5EƐA�~�Vp7�""x��V��j��7�(���W"�A1=���K(�Ѫ��n��SR�����7����?}���=�qR���J'N�cai�K)�m��F��D|`7���C=�in�1�y�-�%È�Q!Pq60�p'N?�b�$r��!�_��?������o}��#����l�g2U�7]�^ʼc%SI�#��\XI5TVW�J.&P	Gbҏ��N!�y�N~�|hHV)"�Z�l&�.�E�Z7nn^�xa�A
2�Hbxt�]=��#p{B�68���PZ�{�$Io"RE������H��ؔb>-4K7�Nk�����?� ���
%���Ӭe��X��JY7EU��%+2*t��fE04د6MK�Ӥ��XYR\��16�S�4m����G���F(эh��c�p��E�g+*R�l��5�=%-�D��*ayq~ӗBPg!�#�Cx�[oy˿7�f�������_�5&&&L��E�k���-s'�gW�bLu�CDդ�?��'����������*���i6��I1moo7�1Yy�ܽ}CC��6����}��cO��6�%Sb[�Wg��2?����K�jk
H�Y�.��8����M�ڤY��i��7ZF"(��� 'ܪ���������M�~'��eBgަ��I3c��J���̚r��'Ua�6|.�� 槯KLʱw~��@�� ���'@�uo��L%9<�SS��Ӗ�Fɛ, x����:�5с��T�q{���J����-���F��
��~��&[o���P\/�Ή?h5bL^�&��z��l�
�&/V��V���4��>���`n~��w�V��S^��r�$i0נTl1-O��50M�yi���֨�wP!�Pk�a1b1Ӓ����4��ı� H������H�קt�����ҙ����>�m	�z���|^?<(�2�dғ�5�B����Y��/��а^�P^ba�Q!Ic�����Y��Eɏ�fr�����6[+@�j��,&
�źSC��;�\�n�/pO�s�����~7cFd�f�=j�Y%�YF���`��߷�|BQ�?f�Qd8�N�݃{�ܭ�'�$CÄz�k�yk����Cwu�J��hZ��J�g[����X$�Z����!nL\:�չK8��
�З���ސ���@7��q����?:�F�+��^�cT,א�60�����jm'r�&�O��܇ޡ=h9��6�Ie@���DOW��;5u:5s'Ϝ@�-*m�<���}������;P��(ێ_��O�s9]MF�;Pk���nazv��YiVjjU3�.��(���~9E3=y��%�)Tr)�+N�;�%�R��#r�$����@��N�ثd�r�#�2EKp{�+���菂)aNJ�UQ�Fj�,�~�b��H��x�V�K���� �J����2F��wm��}$bq�y6��"����6�6,�}'��V �8鱲�A��_�������,��:�Z�o'yZ�у���P�g��0���p�e5�Mjdt@�m�x��Ue�>3��D�\�&F���r*$#�2|2ɣ6Ģ�Y�0����M���m��m?��bL��F��}�҆h�XXY-�jzܸ�#���G(�
�}������x�i�a�'�Q�(ŘL����J�MW��bTl���RK��?��$���;ob#����&��X���@��\W;�.���V����![J���bfl7OZ��NN���ƠL�]HA�0Sh�	����9�j�QS�^'(g�b�؏e��uR�^G�
=:)6o���=�ږ-�?Q�͎֏�����[φ�'�:��|�Q6���5kt�AV[D��ٶ�vf�}�(7L�5*�&=R�f?�*|��L�M��ya�`l1�v;�"q$Y[Dmp6PQ!m1J|���l�x�jð4d���"1�f��k�����7��*d�N1*[@��j���5�����HФx���H�Ø���)G�.9h�O��s����S��7�l&�H8�g�i�+˲࡭�zUg��#N�ȃ�<ö��0)6��r��ML{#P� )�m��I4��btE���<)��Z枌'�2�8<A��uƖӯ�x�
Ec; ��X�Ri�ƚ$5jTT�qe8�K~K�K��d�Z����"�f9��C�G��>�������v��> ����&&���i��(�U+�����㈄��+XZ_���!���E�BNxQ��s���e/�>r;���}���Q�&�e���E-�z����SGN��^\���U��	;�nF$9�\�9~|���tЗ���#1�����k�p��iTUx�^�~\�jz�h�o?���~�����+�2�^����ZL����<    IDAT�F��)�զ��:�RXY���	��ju��Ղ4�r�sX[����54�y8t��(u��ό�=#�4��㔳�+p��p�D����Q��_��s+ȕp����BJW��j1�=���r3�f6D͓-���p>�F\Ŷ��&��C�"1m)�Rz	�r�3mY,����pD�
7�D8�dW~�Sn��4h7 ;�JQ�é(_0�קN��܍��4�S���fNCq��t�%��	!�Z�b[Q|�~(�
G��a�A�7��juy�Э�K�1*��>�
?Xq*ߌ��}i����aL��goh���UT���J���/Q��e2���~�#�j����n���w�=}�c�c�=!
���9T���N�6�TVk`1D�r�@P1�=�}j�ps�<2�S���O��6/7t�ק�K�`r���I���|X �̼�P��v�8}��t*b8����q2%<�	�;-��S�E�L���ܬ|6��rd�kZ�xk�g����y�8�O�to?����f򊯰�z���	�8��ٵ퇊��U9����z������nsme�MJ��՚S��I���SX�誩4�R�څ����4���_�+v�ц�
E�DxdTx��%I�e�a�9]�x�#L1�X^��N8<>��R�L8�-�x4!
R�?����Ĵԫ��!��F�MF%"��b6���������(	,��KP+�˰�\�j�h�ߢ�P_@.�nO@�
!�%A�%���ϡ	!�J���4j>�5��\b�m�~�bU�^6X1L��C�j3*^�gƞS����CՒ���9�5Ŗ�,�=d��M"پN*��5�F6X�Ψ���X)�fJ�C!
�8	���0f��P�;���K�{d?�*]p�Cp9�ڻ\,�:L2Oi0��_B�Y��Z0ָp��.�+�B�1Z�
H~��Dfy��+8���;��KgѨ0p�������v�/6�S*��{���t_x�x�+^���S�d�H�8�N�Oan� w�������9}(U)�n���C*�^W��Ǚs�Qi���{�Apt�齣�������w���Z�˺|o[͔cv9�H��TsHL;;����u���k�����kj+�d��1u�,�&��hQxUG$Ⱦ;��3��(��&)>�w�s����D���#����R;���o�ν7!Snc=SF�ʱ���p+T��Rc;��\f�BN���!`Q��*&SY�؉��k(�S?��
���J����RŜ�EVR��zP{��Bh�~K��h?jg�@(dĩ�;F��{��f�Vt8�t�1�/�����f��͋�n�㩴J��n7�	RȦŨغ2��"����o�Y���Q����&j,.,+��+_��4*&Y��:�j	��aǇ��Pl��G���Q\O�:(��u���n��~���tO�Q��+�
�ۏ݆dwLN�G�ފF��}{H����$ɨ�ӷ�E��\���Fe&BLB7-�y�ɠ�n����+칼^$�{p��7K�K�B���784�{��g�2��d����@P@�����_הׇ���i)��)+m�������b�1{���H��qk���	YM�� �M�^�f�cZ��M�G�,fʍ�X�PP�ɜ�w��:����� ��z-ݓm����W��ŬPGe��-`��6�bR�	V��u�I�7�O@��o�s&Ӵ��RLK*�"c>��b�UN��	��#���Q�$�����9Ou:h�73}�Y�g��c����F<m�/	T����a�/ `V,�T�.M�����O�B���L����ɥ���KE�2�F���`?��u+�s���r��+1�:s���k�t,�{�к���5�v��C7��������]hX�V<�5a��D�5�ows��ĴFM�ﭩ;-|{�繞u~n�e��+Lϴ��.�dR��kN��̭(J���t*�̀)+�NY5ؙC�7?�PLj�i��t�W�c�hv���R�L!n2om�J��� ����m7�!t�	��}>|	� �;�m��p��hbu��.>�r@3Ǌp��ڍ���7؃|��j��߇r���߁������y+x�K��poW.�Bv=��t&_ȇێފ��E����B>�`Ќ�������ϼ�5XZY���k��ڸp�2N����3+�7;p;�ފ�?�B�jQ���D�@"������s8}��~�7�Ǔ�S�������7����\�){���V��wv9=��� ֳ\�2���"ڼ9nf��u��h�Qͯ���XY���YG�^D8��l�؎a�	�s!E�!�$���>��e/F���Ï<�G}�����*��|��v���:jjMb����C/���ʥ��u�uU�T�)�
%���P:������nU�(�Qʭ5�|5�-���e�-Kp:Ӳ�Dꐁj<ع�I��1mV-�H�r�=�ݍ��5��/�n4"Rzr8���]X�9:�����e�o�*�F��ޟ~�����f�-X�g�9�*̙9y�SRmU����7��c;��٠͈���ޚ�`Ɛ�c����3r�C`���X��Yk��7r��%��F��&[Y��BZn�<��tX��������O���M����+�r4Y>/"ԸA������2��_9)�A���x�+^���J�P�7���E9��7D��Z.Ⱥ:%�� �}�����
]���d��zSl���]^&	Ӓ�h�>�,�7V��ZP��%���������e�tNk������`4�t:+݊�q��2LA�=���[V������#�����l��>�lZ>)<���X^ j6,�t,M3~+ɼ�z�.��E��K T�%L��؊c%��X��XB���Ԛu+C��^bm����XK^�I�`=ұ�Y?�w�k��Pk�X.7�<f�p4�w#@�BAB�R�L�7�{{4���OuL��v���K_�Bl�-�¹S��>)��x4��Ω-`B`� �J--���u~�;�#�&���cO
�Hps{v�� �ه�"�j�P�+�Hz���ڣ�6H���s��>�XY-�A���g~��[7�q�"c�gtQ|�	��'0���^f�mi�������"i���wR[��R6`�=g.����l��l]JG�Nv��2�������G�C@�p�� B�j��<!�Z.Ы���|��I �]�#�/G��SF����A�D�.ʜLE���VN� �����_� 6�!���3�g���KG"�^p/����O=���EL�5N�y�=(�*�69�J����<q���Ul��v�;_O�j>Y�G���
�4�%\?���*����}�����ܛ|~[?�|�^���j����/�G}�ATZn��\�:�T��G~�TKeD�.���N�ǵ'Pϯ"�mK�\��q��^�u� E��~�z=����J�y�w�����ˋ����Ϡ�pc)S��R���pGzPo���b��L�Yrz�S��ڢz}<�����Eo�Շt�Ꚃ?V8l�ILK�Jj�<}T*p�.z�`&���+!�:�RéV==hv��
���|���L��3�2�3�q��a~m)�֑x�}�qU�4=\�5D|n��#(�*���"QnZt��5eml�0�Q}�BQf�P��3���f�@�5�lPv[I> �(��������;)
�����m�"J�W
�0����2��d[�o����w�VG�Z[a*k��%+p3}�7�3�&����j[5MV�9z찅cޢI"��}�w����G�67���!1Ok�z0���\Ϝ<���i�����q�Uލ���4
�%���}z��	�t��{�Y�����Z��֕k��:$�B�(���;:g�$���U�e�Z�
�w��w�]��5�W3Ԏ� Lѥ����He�j_����Ԇм�I��ިʷ�}�l�b��������9���ؠ����6p=�1�K���C1�ӌs/aug0a"�k�o�n��կGt���o��5��dE"��"V	 |bT�F���n�Q���֫Ê��[�V��Lf�T�'?Fd� �'f�� �T�蠶�
�N8�A�^@�T�ωvu��A����Ŭb=n��^�S���t�� KO|'�^���nmc]�,�3��]w߁;��pH�6_���	%l������S\Lm\�R�0\ӎ�c,f�bT�6�
���0 v�ɖ��j�@o43O��,o��6pپ�����_�M�Q�5<<�����A�W�w��9�|�|�|���z���N4[z�srԣ�u����N�j�s��J4L0c���C
r�u@)�m�k�2Z���>8B��ݏP�0�(ܞ \ � |�:��N?�m�s�ҙ %��&�{pEѻ�6�=x��Ҝy�YRŃn��KX�~��t��;b��YD�nT#QM�U��"�ۃg�:)9��}�4�}�RQب�G#:҅
�2?q3�9��m��8x�^D�w��IF�e�6���]F�GP�ǩS'pujB4��8Nڨd���������y֨L��1t¯ϔZ�31���&7ն�<p�@%U�E/}:�nG���٫��r��Y�=M<M��ݴ���_�fcaa�tVT8[#kK��.ٽ{7^���bl�G��T�]��?_��.^G��E�k��5��&=Yh�̓���4MJayi΄���R&0Ntf�^ﰇ��D�U�c0S?�RF@�ZL�ɉ��,:b-���E�N�.�Ã�b⦺�JmfՈ
n�4V�6� ��d03���Ӎ={ [.��ܼ�,�C�1U�>�jUճ�OK<@�@eeI��!��L%���7#L3c��F��T���7$A��=�֏�����xVe��r6��
�����lI�@�nO�������@��=���x�S\ƃ.�'�*"�L�Flg���>��o��-`��GB���=`����Mj��)�hgj|HZ��ׇ�G�	X���'�	n�l���������j�
ت�8R�a��"&VS��Iq��ŋ| /\��?�
����Q#�����5�1<�#��R1��/���J� �cN����� ^��/�|�SݽK@�#ϋ��v��_Xc���z*����h�Š2#H������m���m
߾���V��kP��c�N�4�r��X~��L�5hĠK��sk%�
��A�"�b/yɋ��}@��?�Y|���M�o�PnWPԼ��^f���X��أ�Z�w��i0�{��+�l�p���g1a���>[Ӷ�G��Ic�V1�n�@%�*F�	��.��fR���摹���۝�n��^|?Ν=����Z[B_O7z�qLMN��;1e��B��&���s���q���`�K�8��)]�+�M�����ܬ@;G�����\�M&h����n/>�~`�Gl�6����y����bS����s���͎�#r�}ы^(�M�ҕ����Ї>��W�=k�����&���`��P!@��K~1���5�2�J�5�H������w�E��
�eI��8���_���w�	T�8�>�M�����Zx�{�rnh������2c�3�q�?���GQj8�+�=$�������>�]~���^���������t���t�����g����n�\:#��R�`~a�HP-0~��Ϝ��B
�\�@?v8���^9YF�	�?��UE��B�Y���qerB^_:g��H��>���}�����˨��w"W����Ǯͮ�u�zQm��) ��Yg���rA�ʸx�I,N] jiD|M8[%tE|xݫ/zѽ��w����^l���TF��TX5�u��}�]ىH̃��<���GPn�pqj	3+9t�C�{�3U��n�4�*j��^�aeq�jIV���4̑N�ߴ:\n9�J!F��U)R�hT��*�Ya�L���X�����J��`mm]=ݛS�8�T���:��Y�XC�����(VRi\���	{��O�����ǔ�� ��&P��*^��iM�	��?Zm摐�f�M��0<�C��<<��X#��
�N��m��ښ�1#��AfS���m��b�Ȭ���mS��eA��L���As�q
��b��^�CcѸ�'��ȲP�S(c6^#ڬK�d�hm!�m�Ζ�*�go/"�?���������up�2e�%a�d�o�	PxP���'�ǜZ�z�Ӕ� ����%rdpb�RG��.���z�8�o�'�Z]F8�s<H��8ѝ�cnnFm��������I�����U.��ŋ�O��-�������͛A��X�ŇN�=��`�$72)6P��u`m�	2j3F��2K8i$���j��]{[i�v��H�Ef]�C
ߤ�,���+^�2�������?��?ş}��cNv��T�k����}N<*794⾶���)�|ͼ/�l�8��V�{<�H�{�Q�a���ӭ! �?�+��s��P�1��<��^3YB{u�-�ʿ�Σ���-��|�3S�!E�~���`~nF�n��^Q7��H���}-����J���{��t�O��C�r��I���b�x�"K��iCԚ�m��6�0�� z��O����N��,���ύ�ʍ��-�k�c@�=��z�
-�)d�.]���������^Y�,����<n?
�|��s�ѾH�trN�R�mU��0��AeޚQu�k�U�3 ���,m�@��':���Pr._ͶnN.s�nP���c}y��2����gb {C��~�*-���W�s��]�Bn�
F{�Jzr6�n�D����4�σl!f��YD�w��b����S�������?<� ����O����il,���ٍCG�G�o��1�dW�/B<�6���8q�8&9*oM��%��L����g>�ݹ'9#}���?棲��	U����fk�?1��� ?re'.]��*SM��⽜]ũ����4<(�7�FW�F���/H���=��B��h���R1��*�9�ۓLʚ��tim��hQ��A��\_��VR����+I�F���K/�]��l ��.�P��rc
��h:\(3|���I�'2'M8�U�
*�jNzZ��A����w����f��|�^
`}� �<�p(�cw�͇oR����8u�.\��J�)��p�H$�1~m˩�6X�j�m�з�)7B2*),��X^Z�B�TLX�%��:���=r��f�:�w�حϦ�i�ο�A�ƍ�v`b��9nV�z��Ȯ�u X�e{���:�ciX���w����eR!T+��fʵ�M3y!V�M��B7F>��*>�{:P�]����ͨ��Z�`H�:+�'N���p����>*��ЈY�x���d��+Z��f$j�$�Q�59S[��]���_��X4�ߏl���'NT+���1��'�k
�]�2���H�#8w��ܑz�C�/�����E���_n#�3g���G~�l>����b���-�nT��q��ӤBoi��o4���2Һ�P�`
Tl}�/��?�����݈Ry	�:8�&�^�D��GGS���w���?�a�U|�_����ϰ����c�T�q�4d��6�e��ᴗ9��hRk��wq�����!S�c����L ��>+N��M:[����dei#�;��0@�Ҩ��N�
2*l��i�v�Q��^���>.�?�v��h$ ��ٙ��LMLNJsF��Ç��?�*��o�hWca�e�9y�\W���'�T���̴��0�$7�$�M�[�,oit�gy���TL�� S���3�%����۾�~PQ�����=c���[�җ�TCOOR-C�����&���k)�7����*�����TZ7�j7s��QتO��ұpʇ��edLA)0�=����Y�5Q�;�����wÓV�'ֻS@�V3>C��hW��hU�X�����,��87�Ȯ�ر� Z� ����&��O��vy�g�k���c���p`�N�;.E���#a,�/ˁ;�IkT ���`x`��s�4X,X��𖷽�^ş��_���*6V+����#�!�?�<� ͺZL=Q7zb>D}M��:yӳ3,��k�� 5:���O}�=�{p�y*��@3\~Y*R�    IDAT����B� S#�M/��L.by9������2?�Kg�B�����Gõ};qǑ��177�Ƀdߠ��(bO�������$���Lz�w�a`hXfU+�2�j� ��r������|��hMW����Ja��E��W��<�v����޾!��6Z(�z9���e{����W
�Ԣr��h��I%2*4V#�b?�Z�����.���G�C�Ƀ㞻_ ���y<�����#?���,|�(<�Fw�����7�[V�]hi��cD$]BW0�X�+/���;hl���bT�P��R+��#u@�fb�s�!�`cc���u��M#B����?�e�o2	�urh�G��e�����m��>��WX7�T]Y�*O�9�N��T&8�h��{���p���o���J�����(����1�K?�hö!�%��8+�{���cj[�P�Q� �V�^hx��)]~�MYc@�����O��^/ሄ�����x��G5�Ã��"��P����@/z�T�ѝ�
�,��blǐ�O=��B�^x����O};����k+��xY�����Y:/�l1*�O��V�R��Y��ϥ-P�͠�>��}4��NR�'�xul[�h�A+)V�����0�i������.,����/y�臕��/�����y�t�V�+d�_f".Z�D��U�j�Z�Ɠ! ��F�H��S\*"�L��a[P��4u��h ��pJ�P6PQ��'���d��[�|���ɭ��w��o�<���G?�>3-���N<��	��=}�������׼��K�(O���Q+�@����)�z�*�����@�x���RJ�C��<�Lz�Vv׫�H���8����B�$����5�b.�����:%�e����Թ@��
6	R�V��Tr̞����0�-!u�mM�8=F$K�2|>��=J�XR 4���_��>�!6�C3�B��&�@ �����(�G�"ֳ�*z?�͠Qg����hԲ(��©�8�w ���F�9x�q��i����<�� ?@����-{z0��������S��Y��x�.]���ߡ?��J�{��Mؿw� ���,^����������b��\щhr?v<�p��e��F,�H'�c^�;�]-�\������x��A ��y�{�o|�����/P����۱�C�����҇��W��P��19�*�B���r�RHcm�:&�O�]I��."qc�7���.��F�H㜑���fK5�C�@Ξ=�d��\,��I`��4�C�܊�ˋ�s�(�}�{;�RU\�X��Z͎�Ma6A1MA�I,�NI��G�X<���a��14T�W�q5��gWQ$�R/�д��c*�u�cȤ6��019�cώA��!��j#�`xpH��}���.��ɳ�YXB:_���n�Z����U��)�&o�*9�٩���J"�G.����q�t��I�37U����U ��X���-��۹Gf�M&��b��Rn�6��7y�(o�lm�b�U��@��b:���}ӲY~�@�E����a`s�4�9j+�U��h���T���Δ$�ݖHT�LW���=�����y*t�Q�_&Gư�H��@�DɷZj)h�#�h��ɖ�
Ǆɨ���C7=D��[��O<y\�4�2yB�:�F��%1���{p���,�"�w#�aui7<�H8��'O(����^���̧��?`�m,-.�
=N�ŵ�),,/IT����٣7����@�b�J�fN6�������U�Yoe��`�(�%��;�hy��F�x���sd��4Z�8"� Vp۱[�}D��_�������`�ތl��t� _ ���l���Nz�1�)��.�Db��ObN>5�hn:���U%S;ȟ�b�5���%��J��#��
Ŵ- ؕ��2��8~-#�x�s�>w��YiTx_�zb���;s#�h�������>�^o��vU�j��]��
��5,,-�#�5�}����"������yc�g����j�����t��~.P�^����~��������'���Gpu��>tt��_*6��y��1��#[�*\c^�t��V|.y��M�q*����;4�*"���f�ݒ������㏣�I��C09_�n�6X$0̢�Q��Z�W��Q�9�����b���U�9�D���`���:���c�ˇ��܄�{���:y'Μ�����La���]����jdh~�_@��ӯ|�+00:�?����#O���
�)"Hߊ}��g�G�ۈ�P��ଧ�sq؄�yԬH���S˫S�����O�{����ʨLt:>�F�6*�O^_N���w#[s�T�`v1����L���<�k�����4�������a����[���Oh�;�;�'�T:�hWB�o��*�x��8r4�q������nBrp'ǯ���9�r烨#�S�"�o�զɔ>W��:.�?��I�d�@���Yu8�a���gh�x7���\G9��v��j�Pʮˤ��#�v��5�5tE#�NƑMo�^e�O}�x��ؿo��}\ɮ\z ���?4�L���~��8~��݂�L��RT����2ih�uJ�B,�EW,���6�WՂ�H�5+4y�6�^�I=πDNQ]�8�kW'嫱g�>\���k��*bZ��پ�����Z�����ͪ���I�D�z�(d���n��5����q&��ߗ�e�
qC�^�!u�:^'��6�Ģ1كsC�-��B��
GY
 c�Ǵ~�.���Ĵt���*�c�n�����T�u3V�� �ͨ�����,f�ZV#�r�HH�J�Z���,n��\[P��df
Ѱ��=���T�u3؎k�%���x��З���s!�ZÁ�{�R:��� ���7���F<�,���׮���������e�_��L�Օ���hZZ#M�P�a�
��)2��f�6+�gY�omMF8mk�L�|���A>j���L��2F;a�+a�H@��������̧�>��_����%,��j"�Zi+�����Of{�X�[�����ƴ-���Y�>d�4h���]@�JG^7�W�b��"��,��j�yzV�@��D �^`Ƶi��@����}ؽsV��7��/م��	S���u���+��{=Ŵ��D��kw�"Uq��y����8s��*�UN(Rhj酌��L�O�XE���&mք�ѴXL䆭M�׉��o���z�>c>gӽ>�ĳܳ^��
����Gp���Μ=���=������@�wj�*iCa��=�����	M����#
kZ0M��!PѨ�\�����Y�T���%����2O��@uGNw@#�vP&�I�RB8���^�m!z^��`���l=�E��Ѯ��.�ay�<܍UD�5t8r�>��g^��~��Z�+k˘_�Ӛ�E�lUq�����2�GĢ��7ލKW�����1���z��@l=��1�� �`"���91����A��D �F0DE�HC�R~mycq��7��+o���ΨLLt|�p�\�����-w�.41���{��ąTN@en�<V������܉7���Cz�����O�?�dw.Z	GeA�>��]��uype|yZ��,!�A8���=ٻӋ�8?1'7@t ���X^����M�UE���S�~��y�Yf"��E���/����A���/�*��(�v�N��*�k�p��pw�(e�����w����1-�=�ߍ�ߏ��^�#q=�;Gwh3�����h"�;�~z����<��)\�|Y��l�̮�ѢI3��C��fl<�x=��Ĵ�U�9�)p� ��C���d�ǎŁ���8mć����P���c��bY���7w�M��h'+��h�Er���ٕ�ζQ���=l������ /y�X�A,R�scﴴ��C��t��leuǟy����)u9�:�w���j�fe-��Jz+5�2������l*�
��d����{�+����%�pme�H̸b2A�h�f��Ѐ�dk�X2	���pH���I���֙I�I"U�DL14Ul�,*���f<�*�z�ЬU��0'��5�{-�������،_��S>�"�f�03;�f��B���[_�V����)!�k��x����66xѴ�}O	����U�?|�b�5����x, $\4�U5E�.Pܕ�K�H1-������n��_�
�����DW��5�R-`��'��K��YBf�Y^-`�"X"�#�>4c#8aD^<��l�)�0��Q�@�#�tn�q��?:w�A��25J���XTN��RP�E���F6	t�B�=�!�$��)]8sZmO�٢�.p:P�/��9�w%
�.]�,��&=��ckOO��di��tj���_+��l��}
�[-cX���� �����&j����i_[������z$�L)N��=�����'&��p4���e|�ķ��/z��<���M���ɛ:�f�܏�,KF��5١��Y�=�����AW� ��}j�1P�g|N�I�s����O���#ԍ�#_l mwuMC��o��\՚<b��,N�-]cowRvk�K���Z�+qz�ծ�'����gO"lc0�G_W /��n\�pF9r��,/JG�V75��o�-MN)C�ٷ?�x�$�9s˙"� ��#ع�f�@	AT��h q�/�F2D<5�]u9�:�Up�<-;V�76&���_y��=���eT��;�@w�t����K���a�^��6�H�rb}-�r6�N���kg�2w	Ag	�}~�moƱ�F��4D��:y�Q${4�˱fn��XT=���R���ƽ���=k�����F	eę\ٷ�"n�-�0 y<���`ci
h5�q^VS�0�݃����@�b�'*�:��d7P!Ò��4�y?\LdT�ז�i�14؋;��8#�o;�w�7�i��z�&C;�J��f�;p�=�$��S�t��-7�Wְ^�j�]L��r0#����c@��ҝ�u3�jtto��7(=y��Q8�*�y�����\�6��"VЛ�)����nŚ�w�����TL��>���c{��_g���JU��+����e#mn�B^����Ȑ,��@M���$Z>����|���w4�>�\���$�2�3��,�Ζ��*�di�-_3�L�LzyzjJ?�7�b����VǴ��3��l�rۿ{7����#�^Go"���y\d4���}^��˷��ת���:���Ղ���gH]wWB���
�����N�����7�~뷰slL�'���O�����V����j��L���j��N���4�[t�GYN��k� ��a�o:���Aȯ���v�����JR��u��ѡ`�ee9@�`��DWL�˩^�?�ܟ�]��/~Q��)��������%?Ȱ�E�2��y�A0�n-�p�ԛ�As�FՌ�k�6j�#}r�ʛm!���*J�:[�P��M�)6Pi�B?f�t+�Ca<���)9Zu�v��8��6/Y�+�Ǖ	d?�dFGG񶷽��˿Ч�M�w��y愮I:���@�c���{��Ph��ڒܗ�6�~�w�̸�Z��օBx#P�l����t㞲�e���X�jdL�����^��0O ����s*?x�Z7�i�k�r�fY��J�sy����	�6j�o3�.oD�rKd�k�cw(h%�_�����L��'> xp��rFQ�7�C��z����v��g����g�25g<?VWL���]�u�8P+�c~�<��%D�,^:8�{a�}�]*f����[�H��ͷ�%}��U�7 r�d���j*��\զ'�?�#;�@��C��a+��`̃D��������.#W.�)g����j~#�mU������G�|~�J��q�l4��V���ZZ��ȱ�r�,0���6r��
�t꘻~	�S��mp����w���h%��.��ķ��0�52ՐNg4���y.�F���߯�f|О~pt�FY��~L�m��|c�*Ti-SB���&'1�����Obz�<��!W0���;����p�w��Sk�Q���W�*��O/��,K�R)椎�4�*�#��r�1t���]�p(|���.�;��"{��������/�)��ɧ���Թ󈄓X��q��-V<�Q̣v�C�Ң8��xЇHЋ|6�\&�x,&�sF(X�����?��7�]��U${�ES��j!�ǉ��?��5^��kj�F aFN����)�CGl��V��eO�l�>�Md���*�j�7>$*|�PH�%{v�)�릛!�a߁}�����*>���7���jW����TՐA"P!�OPa�9�ٟ^�%�B!.73�q�W/���ᡇ����Q.�4�#���%f�I��^�r���gN��}�:z�1\�t_��o�X�l�t4&O��{rs,�A�M�p꧘�ϔ4U��'B��я|��O6)�?|�1U���f��� P��g��d���Y@e{+�l���~���I�놚Vݝ�c�o��Y;���f�l-���q�G悖�;s�4�՝��O֐��s���������g����B'���c�и_�|�S}b�,Ѯ�u�h��J�Ɵ��l�]��/ɀ#
意~��δ[@�Z7g�hl�B����dTB	jT,��`�)襱cC@��}�:ƃD�?�𓧇���w��xӛ�$ݟA��;���O꾯,��GSJM�"��ƀTӒ�k�ӭ�{l�"�
����֏2����[����γ����6&u����L2m+^����>���g����5*���-�	��:2�>�~�ѾfB�Sf|	��2���j	��.i��::N/j:d{5%T(��4�eM�6�y\�n��C��"F���ۅj�^V̌���B"8�	#=c��w���F��E�z��U�Z��tHg�%�:���q��98ZE&CH��
���ֱ[��ev��	�-/���u##m��ҹ<��Sh��j���~{v`��-��A��A��A��γ��Ee͍_�����#��H\�jf�@�7?��w}���Q!P�Z�ޟ��>=����퍣Pw#Wjcfq�JS����:5��M��S�.b�7��y��ط{Ĳ�w��'�i�`.,:M����	��Q��D�A���r���$~��)�O.�����]8�����	�0}�h�풐߁��	iT�g�ȸn.�P$��Q�H��q���F�h�E��%��+(fWT�jŬ�g�B>/zz���ݧ���w�DOWRU.{��Xv��%4KwP*����=t w�y���o�_�:W9Z�S�XcZ�X	���:�
:��saP�r�T�#�skQbR�Nْ"Py�k^�w��;��͸���X�_+��׿��W'������]LkӴ�A��&g�U��$��Q�7��Q�����7C{c/ܞ��e6G��8�[����7�����"HgS���1�������6�@X��	3�<�Q�Tl��*lC�
'�L�� �̉�g6sF���㗯��PLN�#E�� ����X��~����y��7�!}[�lo��ޤ���MV�zNы����a};;Z���=0by��c�M�$?�+����YYYgWuW�w���-t���a36�6�Np�w��̀H�a6&bbcf<�B�@\���Ё$tw�Z}��ufUV��������R�<���B��UYy���{��{��Ϋ���l�p�-���;���{�
��V�blؒ��m��LNYH4|�a�یw��%�K(� '��ٶ��� �2�2�3i���-PQ��3���PP�v�pD�ϥP�BQ�$~�Y�O|���$p�=��k_���#0���>E|�*�q������*y���+��;�b�Y^�&�Z��BcFF��|v�͖@.ݑ-�B�Td��*.�,P�C-����Q�!����ˠZ*�7M/,����z5IES��1�o���e��E����Ь�4R�V��Ԭ" �������ws�LA���5���2 �Zиv���F �F�
N��0�v�f�t�t���E��ѷ����/'+    IDAT�B���_+�uW,`Ϝ9+���~f���cA�*U��bQ�LL�c�����"Cs�q��c[�E���[���#���e�8��t-Q��	��oyb�D���� >���Mn���K�L1��/ls��4��Q���%5ۺi��Xd�9AJV�Y�+�V�'p��s�4�8zp�^N�0Л��n�U&������y;uꜺ�g��9�ɖ��:M�<@$�M�`d�~�#I*m4;A1�a��0��7�B�e�ʩ��ॗ���v��i @P㮯ܵ������8��7̨<��������j���.�v��T��&g���3W�>#m4�E�gp~�$�fN!�k!�*;�0u�۱�!I����M#�Ԟ��@�Z�u4���/�����?���K��?>�ɹ���<8r�P�zQ�uСwۀ����
�42K�(�VЦ~�T:\��l9�B���LQţ+qx�$�JU��Ey�4*-@�@T����WB[�$n��F�	l�4*��K/�ďT���X��qq{�ɧ����������9��Qi�Pt�n�B���T�:��Q��oN˨���b�@���.��\(�uQ��ٿ~�7p����
��nlG�p�bcŔ�p�0)�f������ب����{A�*��(�2��X����ɏ}��`���:W\v	�})�lA���J������}ߌ*�p)��C��D��@�Js<
 Yx��L�Zgc��>�C2��?7+��l|�sz�>$̘q{�9�Nεu'��1ԢΕW]��#~��h��y�m�!����oߧ4T��/������ʰ���q�ݬ�'�Bm�ZvmZΓ�	�g��z���ѓ��ܹ3���fCM��PЈW���K�	h�q`n��]���^�H�2*�������lGڍʀs�qc�7f1��'��g�b����q�t���sMN����3����ZB�" �0	����8�v�C�O��sB�h4���ATIsm�ՐYY6SC�8����A�|~�J��)4�HtkT���6�J�$��b뇛2]�y�3/�^)#�X~	�F�ɨ����
��r}x|x:xo��=�����^��:4���E�&��e5�l��W^Y���~6�o�i��ǫ�Px���m�#/l��>w&c�G@e�ݷ�����=��7s��^>88(F�@��"�N�9����%��{�,@6g�<��>�h���Q�ǒ�eC�� d�V�Eq~�X\��Ӕ\?���#1�EZ�#���b��H�ݩb����4k���α�%��xg}�OX|$Ԫ�Tx��yi�:��l*����N����S�g�{l�Z�#�����q���x���r�0=���B��!n�7����^lޅ�-{��PsQ�B����~b�6��.$#@�SE�]��ǟ�K/�@G�WG���v5{Ѯ���ؿ���9��Q�F�\�)[��q>�=�	��*n��,be�$�t��Y��U�p~�$Μx�F�F����x�E����799�5�|����N��F�Z	����&\z�a�t�y�)�<w����ul�y	v��t�4=-�Ш�լ�$��_��/�T�ը��V�er����zͤgr��RP�WT8�Ӯ��[B�7nC)T�y��r���ݻ��ށ=�v�Z�����k*٫ɀT_f�p~a'N��#�xB&�{�D�R���)4�5.�L|�3͓	��:6�%�P�e��b[?Ծp�ƶi�0�����?������q:֚���tg�L���#`�2�f���~Y@�?ͤ���m�u�g�7�*�?���� ukl�-��}�����cD��^�"�����a�B=42��Zm���O}_�ƽҟP;�͔ ��E~ɍ֙�q��,P�`��/dߞUߋ�1`��'�AzT	�l:�/>���`��'h�T�ЦA���ޥŖ�3�$���O��v�/ڬ��Z9��(���լ���G��ɤ��hHg�FH�:st\x<	b��q\��'��,�?�Fl�m�K��wn�hˠ�asU�sf�ʫ����:�D���uY㼩c$G��z�3�I˄��LU��xSP��w9�. â�L�h|�n�/1!�p���Q!#g��m�t��)��<":f#����6�m�5I����C.�y�!:����[36	T:��#��*��B�b��E1�l���L�RX[����P_B@��Դ>w46�y�{w�ؔ��_*��ؑ��DSjY�LLL��m��h=(�q�f��޷vP��a�WN�[?�@���uqtw�pa!��R1�5���|�d�L��iY������$�W> �PX�i�^Y�n>�-��8v@��5�_��Ir���w ����Hޥ=bzzF�.W mO�H?<�~�B}%7#�7"�JQ�[Fx�"��*��V�����7y5���3� �Em`2t�-�k9��2�QZ��Y����޽�����!���=Z]��xdnڀ/�pr��v`p�.��}��ڨ�<���h0�A$�F,�Bo�������5;�,����X4�iճ�7|�S�����M��Q	N�߸V�|azi�?:$�jÇ��"�Y�!�wK�27y
���
��9�-��:���$<%u)���J��D�����Q�r��������i�������C���̠����7"ѷK�Ut<>��c5J�g�5n�+p����.���t��0\N���I����R� �Z|?���a�����ĐYMKܘJ���(U�ipo������0���+��?$D:{~���)ep���s�"���cfqQ����ԨX��V��8� r�U"�J^�9h�:����;���
ˁV��j�����)|�[�id���rNu�On�y���n^�^���4�8�`�����糀�hf�3'
 &Ȏ@�^*���=��V{��Cj���\���O߾��j�����P*� tV�댊���&T�`E��#u\vIy��+�+ڴ<~��Q_�K�ٓ�G����C}}r�:{��w�OM�ԙsX�e�m7[R4���F�B0(�_�J�j�C>$Qd��X���"�c����ۿ�ǉ
S�`z�ÛF16�M��<��1��S_�y��Twϴ�6e�d��k��������J��L���K��Zi�ƃ@�)�l�XY^R���l}������\gj�xy<���O��(�6���P�%f�������ұJƢ�44�T�_�jq�](��XZ&�Q�&Q?| ,'�h��&C0	��Q��(�Zzv��F�&i����A�d,�z��v���T�p �g���k�W0,�b�!�������0#H<�;w�D������]��Vܬ����T#��b�֧��ꈕ-[&oQ�Tx��zp��.��86`�<�Oki��mT��l"�S~�mZ�I5��8��s��s��d �y^N��ڋGcƨ�R�q2����Ő%�T�Pj�H�bbb��;^x�1$����O��O*5�M�Pi�(�U����I�6��
�e���Q�����9M�p�!��-21��
m���h��v����,�+X]�C���`�gO�V^5Bt�N?���ƒh�:��`p�6$������B���G�D��[Ѕޘ��Q~�Zu<�³�Y�CE�����g��{���O��gn�M3**��ҵ�Z�Ή�̥�� �U7� ƧӘ�]P�f=Җg'0{�f'N�����Pȣ���GĦ�a	O�X�(�qI��|��TN����������.��X�Ց-{��+�i� �M?:���]�	V�U���f����� ����τ�q⤃��(�o��A B�B�J1m���v��&G[t���7%
p�k�����Y�ѡQ9rD��T�ӎ���s�?�|�,,�b%�Co�0��^��=JN�����țJY ༽�zY�
��)�ZYZ���Y��*TNT�����~>����8I��p�R����c'q�=�bf�<jպ/�-ش�v�O�x�[�`6z���ܘt#(�y���q�uhW�8�PY�p�����=ى���q�����J�H�wn�x&5*dTXm��'�-����	��q��иZm�C���g�]q^�JF�Y�6Ǔ���ݬV����7���<��3j�ђ_�'���i#2���T�z�غm��I9���EJ�^m�5�]n��m�f�U��iT�@$@���6czq�3�Ij�ud��y��pƁ����*xܲk��mA�� �Ԩ8��v��q�z���[��a�6��(�0�c�.���N��ÿ��J�֔�q�0�Z��^1�}~�y̽�M� ;�D����?�V���m:����>3�Tl��N���tU�dD��ډ���`hh�X��R�(�(��R�9R^m�~I���[��J�B����(��M ��������x���ȣ��o��G�'��e��-�����¶ҸQ�5��+�_�8l��i��&貌�=��|��'+�h�i�jA����'��w)RT�)ZP��&{��)�b�G�Y�L�)�ԉ�0�J�$���񱼧d,��:�F(�$)����`K�B��`�����8Mϵ!C���e�!�N���8u1��̚�J ܃Ԧ
�eZrrh;�y�ERp�{�� 3%wc�oN��r]�BK�=^�^�aPYP��t:|S���+�(7���s�u�W��e7=>�6%
M�4y�1%��n�@$�Boj��!����#S����������@��PT�zC������h��xꙧ��ɠX���	X�t��[z����|������:�RL{j�xu�����B�ʖ'���J݃��k��^D���G:s�p������Աg�Y�����Wq�L�M%�Gi!�v
=?��.c4��y�P���O����m�mډ]/�?�B��1�7�(=���g��l6��tZ��~'�|�OV!&�fW����ƍ�a���J�*�ZY@Ec���� ���*>�~R�q]t�X��Y�I�qٻ���4V�3��j����㏠P����Z3�&_BU7<�(�L˰ú�~裲��$F���'}�$�
���?Ė�QS�0,�ZP9���*�ӳ
0�ո�d�B�T�-딯3�(�(}�dV�A����%v����ʶ=c�)�9ހ�"tL�m�.�1�e}�صc��$�vn���>
��_	���Q���Pv�Fh��T����M���e���!�#@��W]u�D�Z�0�u����8�*�ՙz`�B8�&wG�>�^w5.>|��s�Z�4��D�j�$S�X��Q,��#D`ۤ��A=.Ԋ9-��kQx���4?���Eh5ƞ>�N8L����M�@9>�}����p�疚����W�L��T�����hc�|c��n4�F���=�֩؞�\�XC9�m�Q���
a�O�Bm�ͤn��~��c��1�Sۖn�� �H�ƌ)���ˇ`(�$g��_��zU�g������o�.lݼ� /�W�����
�|�fװ��V�F�_P�n?4}krj����Z@v��I-4:��{�Qߪ��9v̍�מV�C}����f0��q�0ΞzE��Ȃ�1,�7�V�5)u7�n�-f�O,ޅ���4�)��#.�;�+z~����c	,�z{=P(��;���~7;�T���NP8#�<�,����-��cK�A1��:
a� �H��9�lud6��u@�X\:�b��O�G-��nӴjK�
f����
�D�s�>��>�T����܂lŅP|��-�i�G��ӹ�a�q�6�e�d�!�/A�[���󳨔��d�'+Gc����"��f��P���8D�e�RT�^)�U+�Ѭ��x�G���{R�<2��/.ڼ&i#J�I��f�̐A
���z|��*���3Obj~�zS�Xd|}�Fv����}����go�- *��˕+��֝Ӌ�k���r݃��9L�, _��� 2� X�f�bTf'O��ܜz��AAG��(�cx`�.: ���Ғ�+�H\5�N��+G��B�3_r5�C[d�FT��hAb�&l��*�^1X�fa���s@kc�U�����k�Ѩ�Q�.��_F��C�Z]G C��7���I�V~?C�T65���Y+� ��i�l��PfQ�T�j�����?���9˅W2**��葒�$�"���fTHi�������?�=�����c����S&x���Ź�Jӥ>h~na��O��cl��_X�d�67���e�	���:�P��mٟwӾ�؜1a��bZ?��Y���6&��1e����m��� J�"���Q!P�֦�0��@�^��,�b��X铌�'�(Je-C$��k�L�HD����c�fځ�}&�Ziժ��Kp䢃�`˅� � Gp� Ohs����i����d�"z��J����6՛��ܬZ?���0g�*׌_����'V��fA����cҨ4���EM,&���a��Y�&�\6&�6�n@��j�ڠ��3=����
���M�sÎ(��U����M���o1V�+/��YyR�D4s��O��|��V�->��m�:���!�^/.���r��-DM�̬��n2���i�ؚ�=�O������E&Gm ���U|u�ht�սV���r�T�*h�ܔ����ͣ�L��8���^�$"8���Nh�9����gCȬ��ZA+�+H��45CF������1<�I�_���T8�#W[k��9���`��g<��M6�Sgjm����]���+�_^uA����s>^)���)ʴ(��S�B��	ۚ\�Tb���J�f�&�By	�uo��K%0A�ҭ9&x�:��V�/��-s*΃×\�l����2E���{��kHHۻi�4��EP����J�"o&yC���&0�����a"�|���y4�5�,�GΤ9�߀s���Ƣ�)�$P*D�(7.���3R�&u?~�Fsh��0�m��z�+�����b�ݠ:5�n���%�{jr�}���0����`��h��id����W��n���~:��{|�r�r�~��b�ږ/�z;�bՃ�92*K(��ٓ�w���_���˘�:���sX��Z�7�y���`f�������F)��cq�(X����ǖ]10��F�J>
�|��星N�cbƖR��c�Q$/ꦡ���ZVr���Y-H�D�R)�Ua>CG�R,ʈ+�L�ڟ�� &ě��(���wժZ�<x�5h��ӃX�5����~%rN��@����A /!c�O}u6}�0b� �V�T4��
��0^��NH�����j�1tt�,SS�8}�,x�!iT���Z`�>�������a�SL.�2fKv2�����w+��z �����U�����<n��;Ƴ�B`~F�ױ���::������%f`����D6���~����?�:ߎYӘ��Q�+Km���TL��(�v����d	�+G=�)Q���9�o~��灉�t��U�j�\y���Mo0�Ғ�Rӌl8q�U�
�c�K�8��9��UPq5Q�%���+��6
�3�5{�aqa�"�wG�E�-�C�P[�n�FB�\�&�N��s�?-H5�6f$���c�mH��_�}9��j�9���}}sc�A ���`5FT�E��l6UjW�&��H�d�C����S+���T������ S��1�_Bd��{�|n��FY������'���цG��ן�����;��O���7,����q#�?�2[�]@Eᓁ��Hqy����%�,��b�vo߆}�2+�?-�kj�N�<!�����7�&7Ӫ�C:7�^}�6n�P�P,��d��m���|�Ɇ��)&�����D��mڄ�.(,�©"EZ8O7K�F=��B�B�BF�E#�n��}�#�¡���|�"� r��6�F�	�L$P���\)|.�5�L��h�F���m@S���/,�9��T&��1=s�X���z��B�g�8�����D��T@��W�cd)�f�1�\���24�W9���x��9V"#C�����^@a=���)�N[��dD)�}M�ld��lt���������U�ŧDq�U�h����H����#m�D�    IDAT�U��<��'4�Za@�� �]����g>���]�sd�B��Z��O��<���cN��/[�ֿ4�\����E�Pz���*�g�T�>NЏ��6��UQ.� �Y����E.��f!C%"D�-�; �!��;�`��h���p#�3�`�����#=�W(Tjz�+d*X��O�.��[YY���(W�e�� �*h�$;�u��f51#~}0
(�Ө�P)�i\���H�Mn�m��ڎ*�L��
�����k쑦kN�J�e[S.��Q�/�`qyMz^<@��i�ցJ*P��
o,[aqC����M7݀w���2KbK�m
��������q<��s��r��:�/�����7�]�x�H�(�1Z�g�Z����T�fӴ.f��E�#-��BSW��8M��Mӿ�s8�bdx#�Gq��G�}�NU����}���}]@E��*=�DҶ��:2+�1��{a�oo��k�X��/�\�9)hVl��;��c�E�:�8����׾HX-#�����::�=�vjQ� �Ϸ���@$��)<����}��j��B.�
�� d =�^���󺰼4��̊�ظ � s�7�Te3�����B$���Y�k�W-#R�&1X�P�ؖ�I'��Um����bۖ�����8>��<�n��1�m,.Ϋ�`+���p��t-8Q��D
���h֗�K��FPk��a��)F�-e �q�-7a���صm�Ƣ'&�t����|�E�V�%�]�7��Mj}���,�dThx��# �$s¢�*b�h6.ƊS?&U����sh��zx�o}�-�?��ӧ1??)�����g��~��(���07��4Փ�5��?�٦���{*x<y=m���eT,˩bͱ0��F� ����m��N:57�I��I@�aT4b��Tl��eW�����v'R��JN�_{���.�0���j�|��X*���,������S(:��������~�E�?�&��¿s�Hg���>4�������Z~[�v`׾�ԁl�o����P-o5���\����	�ÐC�l�v(�nK�@�t���ru9������PC&�)0�[���c%������@� 4@˿]~��O6��s�1��
���U���]�9��`FGx��Ҩ$�z���(��#�[ZF� �,��v5�ol軟���q�u;S�y�rf�~$]����r�M��nLή��S������Ǭ� ����ݪbqa��<V�#���f���J;Hȯ��4`"�`=�Mر�F��/�@&[F�����D��2r�R"O�dpÑ�s�ˋȬ�ѨW��EAU�*����&�W%Xj��S�-�^H�V�)9�����FABA/��Eپ�)�4�~"�0'��4bu��Psmt:�]��pl8S��̌Zg�mE�/:�H�&�T��K��Ţ�S�~h����#غm�6G
M)��B��� �h��.<6��n4Dp!PE��oZ��Q6�կ�w�&��b[��v �G��tH�+ϭ4d��}o �TY�8�5<�̟0<>�F���e\��7� �~��k@�T��I���'_#"�h���srzV)bް��DbQT)ޔ'Im�W�����f������P�7�"�^��H�>/�w�U��>��V��ի&��Xw��|}
�?������ Ǘ��C-��������
z{��k%ƀ�-D�'s,;�sa\B9-dX0�e[5w�,��stL�l�핥��d�����d�+�8e��ʴl��B�a������]�=�~��cqi^7ՠƓE���mu���K��Qf���rf�ި����/S�Ẻ�`F���F�{z$R%��;߅��&�яO?�""�>Dzz5	&FE �����U�B ш=�*tFݳc���o�S�|/��"�k���LrvvF�"_*-�	\|�(>�-#������'Ğ�`��]�d�6�6ry칱�X��k�nh�->~+��dt�E�ЂQ{��r���P��(��n�==�)j�g�	#��w���TCL'ϏX�F��I^�h����|��u�n�u����~�]�������'����y���P��r��ꡋ��R�Pm��t#�VE��1t�!�~XĠÐ\�Z���T����E��`�bA�ض@`�F�Z�wr5kϺ	�4�$�\�X��r�m�_gh ���r=��G�ǎ�JMjJi�贍6.��/�F%�m�U	=x�k2��0Zl����]cC߾��?|�u�~�3��#�b�٥��˪!�R�����Qi��Ei�@��thG
N`dQ*d��,j|��8�rU�h�&��;0�p���0�7m���V�
T�.��O�H_��^��z\&��S�ZI}��ڪ�(�eV�Ѩ��l����1{������6��V9�V��f�(������%cj!��X�nj��*�x4������0N��m5���D��Ju�Ex�̸"�S�E�@�G�@���"�QY^ZԆh]�n*�M`�G���ۣ�����"�j
i�bZ je�f�r��sr�0SHܩ�j������3��3��Wl��*������w��[[�Y�
�M���F!��!��`8�L�;��5iQU����[HP�c߹B��xu��l�ju�)ܧE��˶��b�{H9�31J=�&Z'}�����hPP\D���meQ�E!7@��w���e,.�Q*���4��F�9*��utgNG��S�}j�Bqm]��j��[o��ߎ]{����Fne�?�<}�LO�avf�p�k�js*�q�l�a3ˀX�x|Tm;#��L�[��&ٖ��AǀW��<�^k���Ip��n�B.��`�=D8y󖷼����ͬ�;�x��Л�k�Ƥ�fN���Sf�V�=�KtX� ����.Q�yan^�<���~���u��q�$P����Om;���z��~��=(�)��6�4�e���A����ء�Fc�Y�ϭ*����}������O╗_BvmE�^�F177��L�8޳\4���?|7���w�-U-V0;}^�ȉ'RW��IŶ#5R݀�nP<|~{�-[a7O���$[�Lju9�J4L��fxM�sbY�n!}�}����f],�
������PK�x` ���e�'?��/u?���
���ӌQ��i���ˊ_�HP���c�N�]�a1*#����ш�$��3xe|G.���^9}JT�V+�\o˙}v��-��?��?�֣OEA�LV��8�<b\��
�V�1n��RD�j�E�oM���r��f�'��̔rk/a���MQS$��)��[C"��r�d0�Z|<Yz�3ͪ��xh��[�\�h�d2�8�:��"q���#�n �g?�Vu��8X�o���sl��w}��_�b���.$�O��_��s.S8�λ�Y��N�׃j'�r��J�Ӌ(p܉�+�VT��~$�E�[�G���pmV�TvJX[�*��6�C�!	#�
r�Z�&
�Q��Q@�%�Qf�'�y�T�XY]�Zv	�RA�[��������f� Ҳ��jqM@�U��ծ�U����PG�2��V�Qa��V8o V��h�ƶ
ٓ�c%�q|�,N�W���ؘ�P�.�0$q��Yd���-���x�>��m9��;���YA�f5�ٓi"��j��'y�o߾S@E��H �����U1uiV�3Z�XNno�P(����wM��ud�JgH[u1�K� Y~�ɤh��#�-CM�Le.�h������^��z4j�=F�B���O���ZL�TT�:bZ^��`P#�ܬ�Ic�}n���Ki�D֙t��g�D�G#�̬:�on����M*��i�{|�ɧ���/`-W@�V�7�
>�� ��G�ph�n<��#rW&%Kʘi���x�9��G�/~�KؼeT�N~N�?~?���1>>�ɉYiU)�
�R6�gL��v���U���	Z,ش��2h���;s4M��s�j܂bjJ�I�*D���B���!4�?�`�<��̨ 
[	T��ӟ��ۿ�[|�ӟVVXo�O���h$rV2���:��_k�X?Z��X��ޤ�`*���O���FL�Pe�����\�ɩ|������*�����p���U@%6�s,�J��	4bO�=�x,��y;z�A��7��K���K/��������Wk����;n{;��O��X�`�.ే��$cM(�f�Qt(�Ww{��� ���	-ݎU���Q���F�sXV��7�Yp�/�c��5_k�s�|�M��+����
7�����O}
/;��liiY�7�Af����r�
��=F�a1b��К�jj-爰D�A�4NL�����:G?��1̯���e��A=s���-ېY+ �) _j���t�(b=}Gz���{�\6����nV���r�M��дQ獻%A
���}��ɓb+�:�����h�_{�����*��aJ��g"{Pk��C����X�U0J��_,�	Uz���Ħ�jY���`~�ӟbbnNŵ�N���+{�n��s���_�� *�+����������$\*��S�+879�|��Gp~#�ty$��w{�������_	[0\��^���9���Z��j��k����%�Ɠ�Ş>	f.�H��O*o�pį�{5��ln�BN���7�GD�*�,w�*�)��@�bZS�ѐN���D���3�����3r�eA���Sb����Z�r�M�t��Ȉ�2D�4^���~��ZÛ�K���w�ǧd�O�b�]�͠� �Z�� -9���m��5R�\��K����A��$�Mp��]���~DUw+��ѣ݀ò"*��;j�L��Y��B-��$t��|fa�Aq��ؘ���ϢZ*�w�i�^F�79���f\*<(^4|#8㵡���Д���"��`=F�k�7����;ٲX�컟{�i8bF��瀓UԧP0G�BV�ꫮ�?��/��k��c�=&��{���`rz�7#F�Ŝ2b3�"���ܻ�>�SeUq��:6����`�+��X1�릛o�go��)6z�Z�N�����A��&�gP�T5&M��l!���L�RA�lX&�2 ��+��c���{���jUxNmɈs7+���t���5���~�$�z^���9YU��߼�۸�;��2�dq������F�����@�����sE�#`'Ck&�l+������4[\�^>y3s����i04:��|AA��a�H0���:��{���FڨV�Q�4��������z3^z�<��c(���G�7���	Y<��Z�^�p˛���k�zj�Z��^����#?�����;���ѱ�B6Ԋ�-P����\��d[Ԙ*���X ���IQ�%��5��#�`q�V�W^&?*�l����y�_|������:�g�~�A�@3μF���$��ܵj�bI�u��-][��<`�O�7����g'𺋏�^���b^�����R��JV2-O�
�Ujd|@8�/�9{L[��Z	p5�����.Iw(�R�@�1�S��SH�E�L�Kl���Ǻ|�����)���5!�%�������2�G��&�]���
�/����h*�J���nU0<�����/�����~x������+����ܟ}��W�-`T��������S��k{z�w�bs�k8svպ� bc:��en��i4+p��4f�#�@� �L&+�Ѥ�c@��٠Q�[!(/��?��Y��6�ۏr�Y.1/�T��6'\��5��v��^}#4M��3;�6��8��S@~mQB`��dъ��57�)'ba�.-j�i�)�`G��N#�Ƕ8�1cˇ���0=9���	���g��#�I<2���qvz�zK����Tos"J���Nj7�1�����������׌�� ,�J�⨃�vAGضu;���ua#�T|z�u:�r��րu�5��_#v�lUn���5�����Eͼ��4�p��vt*:�|(�֜vk#��27��jҐL0�%��(d1xr��خ!0���3��6������G�"�)yxyq�@ cc[�c�nM�9wN�gNry�J�ԫ����h�)����\�|/=���_�[�;?���O?�QB!����]���pLi��0m�kؿ{��ށ��l�ޤ�T�ż�/=���%�*?|�u�◾��w�^"s���������8{v\yj�:.���Jf�=�Xʋa�9�h�݁h|��]+��ݼt����ݬ��-�b��T,�	L��Bq$M���3�F`�I��������&���=�җ�"�`l��g�)�G�Q�=�r�4E+UV�|�z+S`E̺��@����>�gdX��)�%����iq#
�`J��0ŷN�5HQU��,�Bɘ�ثSs���E!�׽><8���p-��x�Ȥ0�׋���f���gΜ��ضm*W\u%���ߧ��́ۖ-{�E���RZ�8}g�2M%�uե2�aH�P�#���Ͽ5�{դ�s����.�uZ}�U�|!�s!P������dރ*v�T����'?������#=n���)l��m��z�k��>*�`�0�R��V[�O�Q�{E�Q���̤������S��رk7Jk(7<(�ܨ�X�Pi0�`�-�!h�4C5�)nJk�(��jVT��LM�I#�jvX4�đ}g�����I���mN�ǯ�K��.PKȦ��aሼ���P���h�	Y/�A׃DlP�q�C�.�f��[Ω(�ۉ'g&�QW�'X� ��É{n��|�#��^�)��{��������&��T\m_y���V09��l>'�� �7`4&����x�hX�O��r�r͚�ǂ!R�~�=�;
��guC��ɒ�b�Ώj�#�s���)�ba�dV�C��E��]�5�A�(MB�)�������hVK(d�T�h�
����>]#���t2Y�1�W_��۷�ȋ�
���+%U�L}ݱm����x���?��/�Pd���G1=��󙬌���p�*����,"��/PQz��H�p�(�
�q�7�]f��/���VW״��m�.U=C �+��fi=^}uW@V�`�ch��t��n;b�t.���"��v�1ͬ���e��ѩ/r��7�11c�B��]p�g����V4^���I*��t~�F���ł�V�/dV*� �^*ad˘X���q-�\�������P�4��㏙�b�hT��l[jbz����n\~����O~����ޫM����7� ���Ez�<�=I��	zXas�d�@?�v��x��'1~��x�L+f�04܏f��͋�+�~=��cÁ�i�g�ޮִ����?��gb67�b��[f*��y4���-ph�[b���b�|]c�<��n�iz�d���m�k�j,S��s��1��ԟ��f/Q.2���3�d"�)���K�⮻���ƽ��]_��R��!��If���NA}��x!i��t(��|MM���1��-kj�;z]�ޔ������Y,�Qo�ђO��h�	�0`�*���
�=��p�0E�JC��,�B~�m��@�gf��4/Ϥ�Tk++����A�Y��-�F���W�ؑ@�GƔ�q���8{�,�K�x��'eA?�0�,�*����M���J�wk�,`�̫�P\촟+�k��^k#�֩���s��Wk�����*P��l�A{��Ǵ�𼨥-�K)�cƴ��3����foD�I=7p�{�4�������k�+�8y�6���L�����)lێAYcx�%ouWX�Í�A�+�%��F��%S��Рз(���s�+Uѐ?�����z`���\3��V�_랢-ȞӠ��Ӻ���V�S
�2��5�5��5y����rltL~`�&�O;(���3�D}ضuO=��M�C��u����>8��������r��-����|���~�r�ϟ�YzGǛt!Ѓr͍��y�/d��8�g�|Xy�fG�W~&FJ���¢��QN:�i_�M��4�g�����d����� �O�F��MU�ڗ�]LCu��qoj �F�e�,�WT�E��U/6.�5�r�}c�#z΄�	jhI�T��\f	�BƘ��+H�㲲�,-�OG�R��    IDAT��M�_���$�Ә�?��@V��9Jɾ�W\���Y�{�}���B:�î=�pvj��2*u3�M�=t2*^WS@% �4/��T�H�(�_*z=^@�������������9;v�H��b6V�"��n3=���]l��uc3�X���R-x�:�nQ��D��Z�(^��ɍ�B�VpL�L)q���}��{���¤P���i����tzUN`9-C���+z��,�"M�,�;4�7�񍨖K��/�6&Ho���:�P�x�)�Y�(�s��ɰt}@��
�6�`��1<�裸��a���_�'��=$��}e�s�BfJ�����;o�L��ű�A�'����tZ��{��1���7���ǰ��EƆ��F~-���g?��� 'O����Z�����H�z�͛cS�u�,X���N�]@�nH`�������Ժ�v>ϟekĺ�Z���a�ו"�4/�==�-./`�����W��s�����w�g���uu**�hF8�E��Kd�5��U�����g��ڞ[M�#��iᄝۋJ��V�Ҷ�nD���c$A�9~��곈Q�4�&3:F��7n�NT�8����
��O�.����b�8��M���;vl�uo��}�	����c@�BG�՜�_$�t�^���՘vgcሼդu��v��"h��L�]C�`ڞsx�z`�s��f4)� ���]v�4*b�"1(_����C����c�� �p�eY����$�;7F�W��R}bVh���J	;��q~~�Sҡ��ʫ��vi��yoڂD���\�L�厡�0�.&&S�k�%+PQ��l�7F� r�4*%�.����NC$$�[�@[�f-!�5�i�8�rܙ,�:�i���5ޣ�9z/{nT��p�g4�1��}Ps��.��П��Q�4�ġ�xԏͣ�x��015��	�
t���ɻ�����oP9�R۷��}����[[�xB�(7=8}v+�E�L��+/>�Bf	�:��ƅ�YQ��*��w�!zJV����!#��F�����>�h5��8$�'��#�h��)��M�ؼ}j��6UmՊ.XN�H��qQg�߂>�)�%a�*�QqӜ�UP��V}�V}�����Ȧӆ�`�|�0����	��צ=?�������[148���_�?�郘[L#���Z3�kJ���^uc$� ��]XY^Pk�8/��ښ}N5�ض}�T뉋�M#�X^⸧G?\�m o޴�
m��. �Ԭ���`�
p�q���aX��J����Z�����O��~��5Ԛ�+�8ͤʮ�PuD���"9jh��M�7*�7>6��@py9-{sV(VhkҔ�f�� �ɞ+���4*G�6U?��3��7Zx�cF�ɩ�x�B�HĘpQ'���Z�T���	dWWT������>��s�Gq��@W%;kǱ�]۶�t~v���02+i��T�RK��k��Z�w�4Z�N��� >��0?��v����il�`��u���p�QpUZ�H�]�u�놹�A��6���l�^;��������޸�w�f��$��xL� #1v�ى�~��H0�����퟽C�++���@�P��P����V���
�k���n^g�s�#ae�\�kq'+�|��X�z�a4:.�[�Z�hCap=,�/qc5m�.�"�Հ�
ӓ�5 <�4���>L����z�*�g�%`gn�d_����o��{�{Բp.`]O/>�"&�Ǒ]��'�%P�ԏ&�l8������m/�A�(^�bE�VL�mU`�u���bŲh����ݠ䵊n>�
�|�Qa��S?vL���/~���?�H@� �L�
���n�\�y��:��<��R`괶�G`�V(bn~Q�2�>�%�^&j��6mFr`��.�`/h�����Fd�AF<��t�]]��~?�v��T��@T"[2�xhq:̴�	����^c`Ĉ^ �̵ '�B��x�4�1S�tL�;�!пe!��KiFE���6���zࣳ���Vp�Z��ֱA<��O09=!F��'�@��>�%u����W�ݿu�Ʀ��s���1gWk����;ON-���N8@ō�g���N���EneQ:�P�}f�JFf�F�����;7�w��j�7Ul!t�@t�dGV�Z�s��Xn���Xg�w c;"�>?��+�����I��/y�ܦ2\G�3L�TŚ�si��%�E3�h��ة�u#%�a2*d����Jعk�1�]@��5��f�7�EG���K����c<��{�*�&�kE̯T4IC�:�i���e��p���4�q=���beuU�s����7������'&�=����&�cnn�?���x�K�ț���1B�7Aw�c�U��\4-���U8�+v������,�o7;�lk�"|+!d�T`u��ۣ�m�ݻwk4����������7����06��ZMaq��ɨ0����
�y4����l�-�+�عSm;."��� �>sF��\H~��4%�ozẮT�%9�Z*
h0��V��ܚ�2��9�����F�׹��f!�W��8l�H�'o��ʊ�����}��*���~�ع{�:�\��@y���8q��7]Y!M|]2<�d�}��7i��g���e�n�ۺ��F�N��
i���,��:|�X�	��f���J� ?Fz-�q>(��7Џo|��ڸf��%&8����S)ů�������9����t�꟮n����ώm[��5�ug<��1���8��C�~>�}��E�L�M��2S�(ܮF��è8SP�d
U<qrR�]ͺ܇�N�rؼi@6�gO���jڤ#{=�A�ܽ���mN�gH#���_x�y:�03W(av�L�X�"��TN�6�~Y�a�Sw���]�k�eU�!�m��V�Ƶ��kW��My��_/F�ǋ �@��
���'@�X[���_M�l ����4"_�� .��H��y�2E���R�F�v��Q��N��a`p���BG-�(��0N�����I�.�y#?����p/���^^[�%A^SHl��I��c�3��+��}�k|����L�=�b���$�8rƔ�-R[��h�ݬJ�����@�`}t�f����gWTv��#���hS�%ˆB�-����_���~����|�/
T�ejW��/��Z����_B����E,.�aqn
/=�j�;��N�b��1��L�(�XB��i���r沍ւ�,4�y� z���)o�S���űk�a�#�y7"?:|�Z�{��w[���Xc�M�:�.��[j4�����S!��,�����+��T
7��:\�#����j&��m�f'��13�H������/Py�O �aj>��LI1�|���q���R�8�����G�Ȭ,�K��>g�P0d��P�nx��O?���iᢐ�Ykaq!-�����N�rZ�+/dY	�)_�,i�+���d5*��9�\����P7������稻`J3=���,��$�l�"ڟ֑#���߫�2J�������AL�4��=t|�b-�G�\2��dj��b2*���5?#υ���@k6�D<�p4�qb��(��7��p<;$v%��t�+;-8W��n�&�;f�\R�˰4u����q��Q�S8K
�8�x�GgI	�&�x��s�ο�v��)����3g�87��~��Z@K�}s���d"�s�:hs=<�g"`�`��M�k��nƄg��C7�"Q�T�;2?�>.����V`���1���x�|2�۽w���;�m�������;>���u�R�;��d]i�E@&�\�=��ńdYy���MF�n�{v��`��IV�� 8m���\,�)��[�b�s�b��ad��bO�ɶNi���k �K$d�X`0�Uݰ��4�ke�F��l*��22�D<�s�OI�%`O`	k"����G�
�Ã:d[�&^z�E�=3���4^x�j5LLM��Q�W���31[ ��-��}~-@�v^V��m�g7RN^kM��a78�d<X�\w�u����*����}�l[�|�B����<�X�T����ٴR6�m�9&��!�lF�Z��j��r$}aiYYl�����=�z�o�Q����&Q�y�H�H��򾒓�#:���a�x(�H8�lfE��2��D�0�q�V��aw�/ӊ�>l�5�N�F�8!�bN�A*츎0����m�a��ɀp�_����lT+�rxE��
R��zc��c�fnmE�Ѿ�[����&��h�ϣ�|x�oP��w��Y~K�G�G������g
�+���q֫�kbJ8���x�XX��%�d5��H����K��[Ν���V�S�i����+7W.@L���cf��(�X��S���)�\�������E��.^0t-ʷ��o�Z�|hUѦ֥Y5���I�..ʘ�aW{�oÍ�]��;w��������r���ɛ��~��ڿ����~�S<��18|�lg'��|Re�:��^�&M���@%���b!'�ǯ@A���[c��k�����`*m��R�*A%ӓ_~�eU%��[�Xo�8�I��T�iX����m|1l5%v�Y�l�d$� ���en�Hg��h����:����ݻv���ҋE}�� -L����_�A�
U�`�|�DR>+��t���4o�������Vڱx\���~�+�ym0}}���k���8y��N�T�Uc�2!5E5p���[3I��59UF0`�'
�k�A��JZ3jM�0� ǔ�Jaq!�C})�oy]{)be��ǋ�/�_��_��#��|�^|I��ySSSXXX0�U�F���De����<������&�1'�3�$ϝ=��|�~�&���$\�;��TA��(q����1�������`�4��ܵ���iq���}���.LM� �mZ�ίQ-Ҥ��^j �q��:E��6r)��Qk��`�Ȱƕ��s��A�a�5]M��q��Pi��ғH�\o�J��a%!�q��ց
3�"����9�Mc@#G���zY�M۷K�F�"@�NSwu��~��-��?x��c��Mh7:p�\���8��q�<y����'���	�t�g*l3��%F4^o���jV�`���u� �[5�d;l�i����$�+o`�6��e�c���
�Æ��ӧO����w�_,�A��OZ�s
��-ш1�l�6ۿb���v��ƃ�����N0�1w�z�a�Ʉ&�8!9�����l�w��V�jMo/J-�UG�����D�h�V�J�B�/�&^_��7�� �l��-!����RhV�rC��L2N�SC�k�)t���b:{���Z��*Y@��C�����,���5MD�>�TO�vM�B��E>�AO<�ݻ���?����hp�:��|`s��>���o8��7Ϩ�/��j���Vom��hz�(T���΍�
�R�gZDlmP��*�y^����X��H[�!�Nfg��ɢJy�7;XY��m�i{̓HKuR�2�b��d��S���q�^ԤQi�O�,J�^YNB�E��P�Gv�]C�^��O����d�D���e a =�
k�n�������;����Z���$`�Wۂ�a�=���$���C���ǟԴ��혞_�N��\�DK��"U�~8@F%��r	�2�z��`���.:��w�BЏ|�C�`���:�s�[���I�{�}2��W����ǃ7���_��`o�7#����d��ݺ��ܘ���i��id�]���:�`C6�Ё��D�8t�����E�����������-C�'����eMӔ���H�TF�b[>�0�κ|�\t�P��i9�����ˤ㫮�
�R�z�]�L�N ����p ��C�Z�(�5+9;���
p��-� �#�h��_��XM��ݨ$7�{�v��Lc~fR~Q�dIc�ܹo}�m8r�u���x����ȪP�I��j�c�dU���x[�'��Z�}f��yc�4V'��:w�s�;݆aV�`��m��VP7P!�P{V@θ޲��}@��js,��P/�T�c�ǎC._�:⧉W �P l@@��˜,2���ҔN�&[\Nҵ41��5ka��/��=W�0�N;�X�h��t	��3Ų�x�?,��'`��wGDA�D�Jxv!©�`X?$]�n7z�Q��\O8�X�o�V��!!�F-���<n1*7�x~��;�oӱ[^Z�u���Wd����p��^L�L�B���-t��ۅ�5�
bQ����-{�[���ЂovF^M�a�Nƍ�����E����A�i����!�g{��0��:��+Z��c�(�X��*պ'8��q�珙�ʴe�/��SF
i!@&c�1p��g痱m�>��B 1�
�T(6#�V=�ē�(�7���aLy�x,���0BV�#$g��3�/�o�_��j�}��WP,�`ue	�JA��\v�fM��ı8"[����&���M�i�1Wn �/��j��)ܩ}1`�b}����p5+H<ƕRV�ʎ�#��O~��	����q�N����C�ɿ���3�T�h�ؼ���ʛH�� j-/f��8�c�iUN݈N��T2�a԰ё6��'*���I(��LǭT���!�Hv-[B�T��$Mˌ]0o4�nq���Dq�]������v����x^���E�%�d]a���K��u��yiTdT*Y��E1*h֕��@�c�����{ �}�ס��^�W`Xt`�(R)����'+�I��8��gǞ��ز�HV�b�V��~.���I��b��LR"��D Q���z�ֽ��������$�7������-��}�w~�w#���I��{��ފ{�G�K�-���wa��>��/_��s�/��'�����'q��S�|u+����6�C*v|�F%�	��6w�
o8V��	Tzz����{��$=d�\^�D�՘�<���ۯ�:��NV��e%`�,+���U�S�s.��TlE��j'>��d���NzXF��#�S��dY`��f�B�&���uGŪ��������G�$�������>������e|^2%d�_���A.D��.N��G��p,���6b	3I&��Y~v�����a��_zш�ި�p��rᯔ��°��x/}���ŕ���n�n��/�h�~�id.���#��$H���@��5�--*�Ό�B@�ךP󘘜)��1X~7V�ժi�p����$�I>��"�L�؊�Q���z�s�y1=�׃m�-�nu)v�S��q.�f�t��bK�ϱ��&��.4Ʃ����y�uݴپlj�K.>�h�ǀFz��f�Am�fS���$cA�<]��!��S��Dcn<v�|����K��
X���^����)zhx�P �T%a��g,8]���h�i�v���#�+TK�M�5B������u���E>��?�񣇥���C���Ҽ����?`�G��(�us҈t)���i�t#��U�sf�"����:#˲Z�}�/�n��^�qV�f��a����kp"Q�9�˞�o2��z�Dj�-I�B�5���i�W�5��x�4�P9m��e�TM�` �|�\�DRb^����U�Lb���@�5wuw/Z����q)��f���u���e�P�hDl��ֆ�K�%-��RG�Ű��tȋh XY���K��<Ph-U�p�0-f��l��h"ݫ��Ȟ�����)Ր�n��j}L&�F;֠��i��&���m�Of��B.�.?5*l���ϢŖ��������}��T��G7��ߜ]ȼ��A�@����jW�.+���bv@P}P�V`t��pf�]��SC4�Ѫ"!?6זQ�g��t}kK�[(E�TS{d�D#�B�"�<	��-D�)�qU���h3��$pQ���\���6q�F���8���.��:��h�@�]-	����6��'��󢿷}��>'�~w�}n��f	WV�p��oF__���Ϝ��/���sZԒ�r�}��elm�2�� O�Ȼ�t4�t�Fs��*��q��"���������O��������Ѩ�rz��>��/齈�r�I�G`��Z�bo8[�jь���y    IDATE�-0�l�m��j�nL�G���b����v@c���Ɲ�'0�?�c�h���#�Z������~�?���g�9`�}����i�, �&����V���`Y-���5<2�jjaaI@�Y/ã�x��q�W�u<����MA2)+�6[�����Q<����|-��q��bA�L2+�zS�>0ʰ�	�!|r�ƘC1�:�Mzb�2z|��%��X�a4w&5Ks
��C�M�{�oM��L{G� ���[�Nۮn6��jKl��m���v?��x,��@E 7�WR$����1����@�(lk{$z�-�0@��}9U�uL�ˌ�ݥȑ�?9{i�C��Z���D��}���Mш�&�`4&�)���l9F~lװ���l��m��S�3�J����-p�ASJO�G���@�J����N��l hӨV
�O#�N��sz�1�2`P�a��ѥf�SS��y��U�7��7 3<2*}5-Vӆ�8�Y�h��@^���H�˸��tw�^o�}r�æ�k�
��x�\v�Tv;u��5XͫE�n�5-K�5É�9d]�x<P��O�ZA8�^�̌���'9b}W����c��e	Q�9�ql?��9wi�?x��4���A�B�(5i�F�G�j����l+�� LƻT�cEV��/�gf|q��:�w5v��5�Y��K/�����f�~f�p]�k��R
v2J�m][��~<rR��V�_8�`��pk[�ȗ�F�QH�f���>��j�?�t,��v:�q�(5����1|끯���Z���~��Gc��x�����_���BL;���*�~kvi�]*�����k9\�_U�d�"m��Ȏ�x�x;l_l#�S/�,/�*��у��W���_x�@��H����i�E_�0*�&J��x�py#py��a��Sl��dS�BAb)�Cvk]�O�����q�8}SN�8�
�J�\D��Q�QɡU��C�!h��Hd�4_nL�hz�	]0��c�8��6���:�)�K�.a~a	K˫ژ��F���M�`~y��W^��H���R��/P�X�FaIon���l���y(Ԩ:rP�'�3�>;�����_i\� ;@Ŀ��򜱧�{�	����F�.�����Q��_\lUe+oQ����x{#��]�(��P��z�jc���i�9u󍢂	��خ��߇�����B������td=�>�ɳ��X�:�LN뇴�6[%�v��T�9z\,�?{>W���f�Κ�w�����g�?FCas>���Œ�z�|�x���pu��D�duT�Q��f�{�pDcҤ��ر�b,C�Mc���
u�Qɬ�bsc�dA�8�k*�t2!f͞/�ѐ�44~@�N�������A�}~'��
#�����*f�˞W{-�\)#���������T��ڰ� q�s(b&0��eۂFԮ�h�5�&�U6�\ߤ��\�,hv��m
�H(�����h�/E"��DDL�!g����� X��J����"�29�9���s�Q��&\�Dj�����V�l����3̕1���A��hk3�.�x0:2��W�%�$B�5����Qg��l��0�����!�;�@:����9�l&��,��Ҷ����V������bIDo��,���?��,��>A��k�^+����^K��<��6x}���x�]&��o�Z]h1�8dR�	T�M���tk%f�(�CN�5�;�27�EZX��T��Z�p�|����r6�rmC��0:y5�Pu%�	��v�C#d>9V���1ϹK�X�j��H���5S{�)��Ջ2�M�U�`��\{����	��z���TB�'[Sb=����y8�Q�.k|~hd/�!�x��3hyBH��Pn��v)����V���HH�����nqҒ���L��7��U\�F��͉�i��ͣ㽯����������ygןF�c���f�-�R'�Tc�o�����%�V%�rv	Ks�096��n��Ͻ`����w�'�م54;^T9sK"N N`px/������p�	#M��f�YD%Gy	H�yi��r���6�R�K[���65��*���bZ*�iq\+m�Q��{���F�@�c�q�AD#�g(�OFO"�|�X���y���Y�X��V��� <� *�V:^l��A&�������a8�+���RC*R�'����c�;��[&F�}i��oǿ������[pè,.��/�� .��;�X�Y�5*���eTĔqv�aC�x���97	~�g���v���E��m)f-��*�ZF�~��!�n0�ц��@��ԛ5���O����s	����w;@ŧ�n��c�6�6R�%@���J����XB*�������I-�F��fb�@��o�6>&���-�t�<vx��Q*�6���Q�jO=�<Ο?_0���;����-��Y��;�ަ�O8�G<@vk���2�����j3�۴�r����Xüq"����i朙M_>1l��0L $Ϗ�Ͱ��Q��ڴ_ʎA�I�~սVջü�G�e���~@Ľ�2 ̛	j��HL�+�Mtpj6|/���	���zn������-l��F�� h
�#}2�#0`�#����Q�b3}ܠ��.po;]Y���>TZm�kJ��z�fD�n��QI$�]�5�#=��=�K$P'C#��X�3�%�� L���[��HţH�cX]^g[]<teiFM^k�|��t��������� ��V������@ES?\n����+wa���<�|��-d�Qsϳ�lϭ4;k�? l_V�����֏5���z�H�Z����뎠�?׽�
hm%����I?�+�7�Z�B�R�(�y��+��1=\�X�Ɔ1�ct��qM�-��ax�~�LA�A�C'4wx`�T�]M��K����t$I�"�v���T*%�qR�(�Dx��"�[�y�l\yEm�C��4P�����tJE=YX����i?��7�7����M���7̭n�;����Ø�_F�K{D�.�X$�DăT�O�f�M]����er�����a�δ����\�P�x�����_��[���s�?���:���O��O_��|�J�D����j	�g�]f�8�V�X�&hm<]�m���X_��ի�5�S?��G�-�DM�g����1^<{���X�d�R�[��F S��O���#�ZX�,��	��Z� �Pr����R!����T��T��1x2��,�*�w�ꐹ`��Z�
�T�Rrg$���H�\�x|��gF�O������\>�����W� �W�a~q]V�S��|���P1�+7��YF%�Q�n�amuY@E�Ù�go=�����O�ԇ�.���j���������/�왗�o�<(�R��-ñ{!Q+��]��c�v>F?'Ǆ�-���w�,0�7q�u�#w6B�r�B[C�jg���T2{'��v����*ܷB- nF��O��?��?P!~�fA�F2*��qdt�}r�tsdO����"$�7�O�]�� �fe�� �3>΍�q3�6��bo���5Q+���glG���P���]�;-�}�Ν{E��zvp�5U����ۇ�o��l��P̙�g2nZ�=z]ۮ�@����n�U���(�YPYQ-����kU�;�wT�&d��zN[�jv��f���|SH��M��h1yC����$�m���d�8!�m�0F�f�s�C
=.1>��5#g������6j�h^& ����A����� �	����T�5Tj-k�P��P��{0�ſ�	p��$fy���l3+{�:����򨕡@i�NoR�����^�-/�c}kMׯ�j��f�����%��a1*��sڍ��؞�2-�l�L�)S�u�P��>[�L#o�:�g[�Q�����S���E`�1N�p�=og�����^�cF�	2���F(�S����kkԛ�!��k�qx��9��`��7	NM�X��<r�;"��az�%İ�յ5�p�)�nfpmqC��0���8���dKe �&�}���:[�f��SU�(�Z�ƣڣ
�<�����y,��B6�<{W�>�t�������Ǒ��&M���O>�vT���h��'���~��	�����7�_y����c���"9<����=ht��*�Q�����	�}��� �j+x�t��%sӉ=�x����Qi��;%Ǔ�����}�����u�uT�G�֧/ͭ���O������J	��)=���x��0:mN�t�m��0s�g�E����d��'�O��?���D9W+m<��S:��W�4��la+_[�%��x��`r�Q4;>,o�u��u��M��F���tQ.䰙Yբ�gfxȣB��c4�F:��8�E�l};����Z@�jA�b�ع,ŢdT�(�$��
��͕��'��ł�1$����)��4�f���Ռ*��GO`quKk�}r鵭T��P�b�~67�TD{2�SSP��=��?��?��'�� �z���L/^�W��wx����j��?����x-"��of�v��L����X�����Y
׎0�hvK-�w�:^�F�Y��&M�Ȟ�6��	�Q�<u`��@��g���OJ���P/j�g��ԫ�|c�o���EmC�X�/�
O��Ms�]1f��U#�;�#�jI�3�v���!Q�>/�Ţ@s,�$@���F�z,��U|��T�.�k2!s�=��Ay`�t|��<)�&�F��nHtK�~��#��������f#�h�i�<��9�vD�\+�1�Uc��;�WG3 ��T^m�p#0��{��Հ�dA�5��c��]
��E#M�ȞQ��`5�m�vӒ0V�Tқ\����k�튊����P��A!�E�c��޸�VUb辞��G9
J
��fzdS�+V�+WQe��D�mF�zB���%Y��J}�4*p+��ǀ�J�'��ya%�Q�~��r�}�٧T�bۛ��ի�©�`�5'��(�d����6��{�U ���EM��g����863d�9s�:>*+ԩ�GE���&��߻۲�Ű�.�ml�1��k�f����Ͷ��!��n'ݸ6�ڰ��]�t��𓱢8��D�g�?P��pGY��t`�1�<��yk��2��y<?�3�d[m\�������n��ꆦ3�&0~�8�j���^��S�BH ��/2t�<Yk��.��f��D�W��{��q",��b�/�Za��~��s�����a���Qev����E�9�!��ː�7�Դ+�ѡ��0u�0.N����_�f��s��_�b��q���.�J
sl�'�/7�h���h�J�ɹ���R�H CҨ��͢EcA"�W�n���O����̭���F%��O]��xw7�#�BFea��K3�;��p��{S�R���,�� �2�@����}���{�}/���w�ѬH����w��v�*����*r�lך(7(A<݋��<b��M��d��l(UZh2(���g�&��-
��(nTk�	�?i��-	TxrTȨ���M���;�ƅ���6b�X�lfǤ���hY��X�('��ʶ�?-�z<��m��3u�(r�2�.,J ��g��ZQ^ը�'���D �᩹-0��H0 s��o>��������/�/�ڵy�>}/�}���;U-ov�1Y�b{�v���o*���?vDP�#~�Nn6p#Ƴ�����ֱ؉ 3
kl��\�yyb��,
�ET!������<r_��K����#�2	U��Ɠɨp�=~��X1�ދ����1�`�iMt�#��1�^�@�1�;$&���8Jk����T��#�Nk�m��N����������|�\�_�x����V�Պĝ^7�:b�ҡ�"Ǝ�)�\Y_+ �� �r��1��x�n�E�.�Q.[?|L�Pv6$#�d5m�.~��sLVB����q\1-x�����uj6w��lU.�xW[Jt��L���� �4ڈEz���UU�&�ZU4=�$�s����F�l���i��ǆ�*�*�����I0�Ǣ**�[[�3��K0�E2F]��ǰg|�H�JYm�z�.�)���ͣ�1o�OԨ�8IFf%��G�ii^*|�.D���_k������0>��w��z��ob}mѰ�=�_���:�r��#�҉0��Do2%���?�]_�����M��ɩ*�-҉�`X�T��R�D�R�K�T+�������3�i����m[ݚ=�\[&�^��y�y����T�5d�X��$m�����#p��{�[���Y��2�1
�YdF0I�jB5A8<���yH�TZ����=q���XZ�@��^�:.F��|?�~zQ��r�l�0�j&Q& +{S��J��n�50��"��y�S�q�'�1?���&�z1� �f]F���*��e���h#kϑeEt�ػ�:�_?.\����l��ǟ?���-lm7�w�R���_�Dq��@(&C�x��~�����.巐��or�FLK���s����#�?���3����� �̬��m�ݟ�]̼!V!��,�p���
g��nW�v�	���\���D~i���NY���o=�����?�Q�˗f��ʥil����EP��$Z�PT� ���[nC4ч'�~�v ��(�8�D�c���t�9�XZ��F�,�J�P�XRؤ)����㥭_m�Q�@�C��!��^lC���X�<m�!mN����������)��a�b#���V^l���ַ�XX]W��)nkp$���'c�\O��8GoD�*��e���u�8R�s����E���)��4;��֋#ʴ��w��v&[����bM�X�X��\���([Q�h�x�����lv��7����_�1�̫�ʪK��b�;+�Օ5��f�P��'��'�sjj�2>�HG陽B�aFߍ�C���d¡�w�*�
���X#'Qፆ6AM�8c�A�w�54��ڏw�{��GV���104�1�'�y�����N�;Ӯ��94L�vw1ڟ[~\0�P��G��YC6g<FTQ����������ڜ�6�������[*������K�|�@g���*�j���w�:_�VT1;��m";�l+ns�\
��,�붒��	70�l���f�{������d4�#��iz�a|dؾ��c����;d�YD#	M�Z�F�+�*0Þ0K\je�Q���b{��+�bt�dx��RSA#Ky������ra��-��/7�H[(WuM�aj�M�
���aq"1��c4O�&��v�O�Iه���{�y�f����Ocmu	��I�	,���x����n��H$��={�|L�s���h�� �+����c{�`m}Sײ��5� �cu*|�]~�b�}�S��9dxNy��H���5��߈�)~6Š
!��Pr4+�
��_�s]a�����@�,#������y�Cw�o ��H��5H����ף�WO���Z��p��	1Q3W����H��c��5�����߈�K+�<{��{16uuW5w�� ��AԻ��!�e��X*y8�(;S�����K�L��%Oa���	�*�x��"�|��N��F~sI�&5\��꺑ə����2�4��;ߤV8��3�Y;qR]���V68sy�9�;r=�?�FldK���x�$�!��e����YGvsM���F�Ѓ�
�)4�܂�[�88������Ͼ>�ʕ����V�����v�IԺ!T�^�fJ��[A�L�y��!cQ?Z�.��,��E��Co�����A�?���4���ɪr�&��J���ǧ�z�;LN�KC�7܊��t}b_��c��M!W�ލ Wi��60���i�Z�#�Y��m�9$i�u"u� T�:-�(*Ҩ3j�4�YM,u�5��Qi��B��Q�b�@:�D$� D�@3��H��������p�%�(Ujkqz �?���-�fs���Na�<����K��H�+1-��=jU%^��'2'��ʑ�V�ⴇmq���Pef��l��Ʊ�������m%��󇏳�!V�b�,\(��ݞd,P����f�Pʆq%C�E���ZMU�3�_�5E>�hT��.�4�ҡ��vILKS6j��    IDATtXU�V�'���|297j�8���=�/���3ڔ	�fx�b$���ަ���mdr���
Bј�ZvK�Ƨ��_���T��#c���?��������µ��)jv�~���}IF����Q+��@�]Ѩ�����8�<2p���>�7���;��A�i�=��1����e���4�
��͂J��qS`�_����6��aHt���-^w<H��e�Ey�؊ٴ�h�刐k՝�
�{0�*��Pn�<�k+��-�}Q(_.�p��q�گ����׊NP4 ]����TG���d�B���]�b����|>.�Ԉо�;�x�x�H|L$����9���Z]���)u��J%�T<sl�~D�)�����h*���K�h��g���q&S{�����w��������X��U맷'!v$����! �h�侽������'�y���eM�������N�����VV��
���*h�NK��?�8�oޟ��4,��������Xc��c�r4G|xv�ݠ�~'0�?�i����0��3�����znh^ob�ن�2��0\�(¦8��mc�ʸ&+T6�����ø��o���U��W�-��6i'n�	�[9�I�cߑPAuO�� ��*��aT@6��ވ���ϣV, H�Lo}��w��m1����� �t����8�̣L�q��T�F{����`yi���YYY��^A��K���;q�
'������3�O���7��l�gq��5$��M����2��<�x�с���
%�0��R�{1�����L[�
U.Դ߯mL�&>�;���^@e.S?��y�����w)T;AT��D�\]B�T���1'/��:6�fp�GQ�/��.!� �����M7��':N�zt��b[��J(A"գ�Ծ��O��� k��x��o������1�T�����Z�+�F��0���I�z����
ZՒX��.'U���1R�ZHǘ!�n���ji�i�Y���M�nˉ!.4D��bA7	��T2��ǃ��l�9��|���9GNN��fv�=�8Μ��1�T�<A��'1����B^��
�i%�u�^F�YC*��bZ)�5Vj�qȰ�p�`�0��0LN�3�-�ё=ZH�G���H������m�Xz�g��m�F[A�\���F�QÊ�8���m�P�oǌ͚J�B7VS|�����b� �T��[�v�4��E���4�D�Љ�bR1�թ�$�[��1=�676D给��"��	#CF��^,���0�bQ���������0��_���ۇ�~��q����ǿ'_N\02B�����6�a?n��J[�:{���dW�L�'�] �sZ�Y����y���V�ۘ��Ʒ�����f��C�z���]�t=fh!���O��1�{��Fհ5Hd�3�l�7��=�h+sJP���ߕ��E#.^���ZN;��0J�@X^n+�`��8���n�m��G�X���?�}��'�h��W��Ϊ<7J��������N~�Y�`��P���{S1i�b��#��hv|:vԗq�7�+b#�C�^)����M��w�
W��w"�(�Q#�$cJf����c���܋��_�s�<)f�7�B*�=22�������9�ʏ��?���G�����PEͩ�͍����G������l�ǆ(k��BMW�hq��m���ԏ�hb,�b�eMvG,�;�}���
���X֖�Ǳc�d�Ȃ�m_��f������>����*�����bЧ�Q���+nŗ�������Z�L!/oo��������M�c���+X�dq�M7cy}���``l���@�F͛BCh���n��!���}��:�͹K(�^EW�A�]�<�ѩc�����j��Z-AO�q��i�{�)�����/�Av�l)�qZS�+P� ��]���8r�<._�(��v��'%�����x��Yx�q�*-\�����\�;��;��#������u������sSaZ?�bV�ξ�1���k�du95I����qd$����?��_�2*���������BԨ�Pk���^P�i��A*��ȵK/�̳߁�[F�SG*�G:�u�aj�~%����N`�i�2)g�TJ:��tZ��z�����҂�4��g//��o>�X�AT:1��]p�U��NAO�Z	k�װ�ۄ�[��a�ZĨ'�J/Th�Ӕ�����M�T,P�>�ȕ@EQ�����P�&j���(n��V��1���v�͢�������k�|q�`��$�}�tuk���
7wc�Օn�Ӭh�#���@�v��3k�vX.4�a��k7���>ݰ�}ê4F�ǵP4���?�ū�o����:�s۲�n��n�r�L�q��p&�,��1G�VI��]�%�/�wt/U�aU��i��	8���%�iu���2��Q��@ŀ������ҽ�4iDc�\./���d�KtL6SL
�c�:�D09A�r-zt�[o�'�;��Ϝ���9Yk=~��p�&H����|eF-��v����&}��p�]o���<.�?���8�?���Sf{ln����7\�_����7�u��Z�wiW�r�
���U���n��bTxݐ&��i�t�w
����.rgꋏ'@��[@k�,��%�e:�#���A	���Y��9�i��z^�rT8�����!�T<�@�+;�;���k�*�������?�	1*�C����I�0͘����m��:`K�[A��Z��&��I%c�I��7#P5�Uf�	(�BI-�l>/}�yP�u�*tخ5x�z�cD ���"� �h��' ǎ�O������x������e� aqaN�eq�$#�@($!9��'~SS��� 2��(�Y�+�\Ik��ʆڎ��&���!�B��<T�y���
G�F��ՙY�����[��=�������f����>�>�%"�B�3�?��?�w���+�%P�4'�T���ˮ��2:�G�Vk�@���]��M�Uh�h=u�0}eF��n:%�r�ʌ�~�=�J'$�≎��G�A!/�\]��q���!;}h5A#[�@�p�#�x�=��۶��Hȋ�t�=�-l,]�@O'���������^���c�Đ/����jucU�~"G�Z��?����d�E�M�eJ������WQ�����̭�	t������D~->�ɩ�����ޑ�B���`v�ʟ��/���^�ʑb���+���G0�#,�������E�+��߃J~��^�̹��i��=qE����*LV.�Ӆf��N�~���\yc�eB&e��a9:�k�fqi�&��Cr`_���׃�;���[p�M�ծ!p�]�c���Xe�R��M�7����>��1��͎�WY�Մ���u
i�Q/g5��fU�\T����ËM���0zbq�p�q�߃�ƚ*���altXN��dL@���|������'q��Q�d�����^�Z��@�۪�o�� ��!�� �.�42̂���)�E����GĦp��O{g�ؘ���w`7(;Z�߱����w��-=��@����| ��(��vwl��F���1�jbmsC�(#j�"i���{h��C0Ǌ;�H|F��<Ȱ� Pq&�j��V�<_��̘��x2G-Ǚ�/cz抨|���4�
xP����P�.�2؛��3�r���CA�^�r/�9�L!��͌2*�:�#�L�R�~�=o���^z�9	i9�V*�O�D����R>/͟�������͔��u�ʷ���XZZ���9-�E��6̈����+wX'����9��&�l'�t~���j�$�s���/��ئsc�=�/nC�rHq�^�u؛baH��|�l�D��\_�ͷ܀_���=�w��>���s�0��+�z_ ��`:��E��wؾ�@E�z]�EA ��R��B�HDm�H�v�]�*�cDj^ʵ�tJ�z�jUL$F0PUδ�����A�V���dnV��䲛:�E~���Ank��~	�s���;@ejj�|P�^��Ɔ��̣�п�I�?%�!��ҥi��LA��9���f����g3�*��*���66"��~G���T����P�oV�$0�~���)(,`�����8���N������
�22*����?�<��C:\��x;�EF��^�c��T,8"�Y����m�-t7���y�00<�x�3�ΣP�V���f�fg��ƾ#'Qme��M��B��5A��B�U���@i�4�a�JY�h�T*� ��^��=@&_6-�f=��A<��W�]X�h_S}���7�8�f��'{�b'o�#��~��+bת�
��j�2�2��9T�秾�Xn!Wi��/��j�
p�;߇xϐ��W��vx ��t/�9��]��	{�wlH@eaiM�{gB�߭nO����������$����G�Q��^�W�x�ҵ����dT*�֋*�B�`\���.��$
�3p��H�|�K�/ݣ,��t!�r�b��4z��A\�tg^���Q@��Z��~<�~�:�&�㮷�K�*���s����Oa=_A]�Ϯ�H�7�q��s�.^eSiR�K!�?�xjP�D�&�k����i�Զ�T��U)	,��Ð@
i	Tr�Z\ٳ�EC8�w/n;u�Ҕ�fgЛ���Р�{p��Q�O�a��
�x�W�o��&�>�b���W�i�@�_�~�it�=]��!$�AM������(��UJL����(�9�Ka�I-��^� ���؄Dy�|XFE�#��M��fL^�O�]!��;��fi}����A�7;	b�����N�4���3(������%n��č�m���]4B꺔�M�p��B!_�X����cS������@�BRn����|�HTS@���ГmCm�����j��Y����	+���aM)ј��W.^@.��ޡU��YW��EWH:�r\6����6E&������U�D&�����J�bN�-�܂��������+[��Ja[���˫r%6FX��&�(x�X<��";�8��}'׉��hgly�F��5�&7_u%�bkn<o�\�_����	"��C�D�8��B �|���$�Q�8y��G14<�/��U|��������}̑R�1��`lk++�|�|���*��J��D!"�P�y_m����a6O���mQ^7�V��XfG���w]hp2Mw�T��
�k<�V�S��R�{�*�/ pt�0�k�k(��t���Ԯ�-���n`meEB�\A�2�	y_s�����8����R��m���X]�P�g}Ӵ~,�b�
��nF�N머qZs<W|�b[9�����ׅebl�O��3Uh[��=�@׶m��2**��z�^�:%�z����70Y>�� �\~տ��t�jb�I5'#����f��q�ư��x�}|.2�˫J����ƛo�zfW�͡g`��C��CQ��c��FPsE�7 �X�bs��/}����"|�4]a{�q����ӡ����m��!�{��X]:���^�w���:y�}X^\@��B*ًvǃ�W��GW�Q�TB0@�R�Lo 
��܈�{�)5pazs�Ed+]����C�w�"�e��:z� *-�[��*{F�����99�Z��C}��h�~�?����L��&k�^�����c[?dT���*��#Zh�+�x�ɇ��:|��a�m1����_~������^���7�o���E�^[���Z��fc[�X:�R�zӭ���y;�y_��SX/�0��8�re���܅�[��Q���˘~�ytY����2�f�� ��'��G�����݂�Y�Rί�YiW�T@�J��d"�d*������=n���`���D_:���&�="VȊ�&�M����y��G��/}/����ѽX��)V���2�ћ��'Pa�ko<��N�T�%�'��n*�i��i�?�}�p��-�4���H1���5�<��eFl����ײ0�¶@�R�̢�kZQ��i���y{�F�B�~��'L;n����C�+��\D/��Z֨�L�Z����f{!O�
 ��G�X���aGI͗�L�8��v�4
_�$X.�lgВ�!w��}��*hn��e�B$���0�?~O=��|1�|��ܳN{�!�%f:-��I�
ElW���ď��������RV��4s=�>\�6��o�I-����*DNy��/�{�����N�LN��'�xJB�+ӳ��lW��QXlƳ����ⴻ����0X���qZ{�X�£I�"��2V��1���f}��X�=֬d5m���s����a{�/�F4D.����q��o�������Ҩ,��brb��.�������X�V.+��	T�ٔ��b��	N>u�{Ь�6]������ M�i�!�=����]�x�7��3~-LP��°�J��n��5K�̄L��jH��>Am[As��L�J��F�9�������e5oL����x��=���6_�T�K/��f�g#cT-+�R��k1��3�>�|Za�d�,z̔���E
��ZGY^/V�f�n��m�fe����C6���L��d"�{��{��+_#��"S"֓Es�.1*�wN�H3�u���E�B,^s�a!H� ��Ȧr:jf�2���=�khie#��w��ծT"����R��,�]���+�b{�
�m����PcOb����/1���C�Ao�_�.�]~{FR801�w�s�v�mL�p��E1fl�--m��3g\#1N���=�ӇÇ ��dQI�����8}~��\��@��CD$ُ�b5��]�L�ݰY��L�.˨|��o��Q�hU�g��H�O>�����_���ba����k�?�`���O�é��g�e�D� 3p�釀�5�5�F�����=~�kXϬ�ԍ7hb���763U}��⽅d"dƝ#A�z���n�<���m<��,gZ8~�-���AM��6B�Us�r�9̟Q�iyNpLN4g �x/�CB���(�Ɠ��Pͪ�����0*����|hm��)�hy���Ǜ�p��B��������C������Б#�(<��s���_�s/�PYX�D��D��>2&sB����d�60���'sb��'��U���(����#�ӂ��!<���0s�*��^��QmT�]��i���*��l�&��c7��?�����v�Vr�fM�8N��6��"�w�-r��w�%h���bF�G�Oi��D*��90Џ��>��)ǕbU� Y#�~�Ѱz�l!��H�*ېB3�	.j|�'Ԩ�
N�S�2Uun~^�:Y?��Ȧ�қSVnN�5[���~/�ffT�{��̳O��%eOA\�XPt���R���6�C��]鬆{��[��X�3-���<�OMj��g���������Moک�7V����g0;{M>:*�fSŀ>���BM�=w���q��}p{�f��5C1�*g��[%[��O��rr���=�*�������⒀*�4����%�����O�'q�����ۿ�ۘ��G<��h:M�����x$6T���p�⨸F�[M���h6*&U��~ ���ļl�T�+�]h:�8|�Ն��x��-�ª>��1���|t����{z�rȶ�˨��4���}�k-2){d�_ka����t9w���y���~��!]זU��hZ?ۥ�
����o`u=cX�ms�y���)�'�e�m�Z0jYk�@�f�p�+�&H�S��}�㾛}�T����/2����k�Ƶ�w�w��� _��'���G�ǞS_��ɤ0�����J$���0G�)h�.��O6_и�V&�@4����������1<�#{"Ws��Kß�+<����	���(�������sX_��V��6��^ć�������]G�ڂ��S�1qc����,��.�%񮷾�yǛ�i7�����m�������/\�Cm���4N�8.�H�y��� ����� {��.e������a9�f�k�N�>
�}��5k�p�L�㑇����;�F�n����������_��;��6�Wm������}[?�F�W.�o�t.J    IDAT���+�zۍ�MT��H��|���yL�y���$�8�c2��Mªgt�(����mltP�|�����}me�z}�	���8y�q��������n�1=���_XVr�ā��)��wao�Zӧ��,�J5�+��H�0��>��%�F�t�0�S\p^*���0*t�Wy��H�đY[7f��6z{5^H���fFdT4�����0�������V�x�,�����3�a�Ĕ|Vr�0QoA>��l9@e0����Fns]B@�l�y�f3�3-E�7�|Jm�S�n�M}��v�k����ϼ �%���:�l4�r�bZ3�ݛ�nZw7�bo���)��u�td�Q����J\T3G@9�<2CQ���_Ǯ;nB�=̊�S�����ߒ8��
�
�5������V� �,�����M�qw��jH$�
�c�{l-p�:hR�O�yϾ�<|ސ�᫵�{V�Ũ?|�H@�1��R+��1	�n魞�E V��F5�;���%��Ҩ �T��2`�r���*y���,¡���~�W~E�;=��X_^Vˇ�
[k��?�ie�e��x��6qg"��_��峛E��᧺��[����e�aI��Mѹ�Բs^��k"�k#�0*=��a�[J����m���(���33��M���"�Hc}s�䔀
�T��ȼ�5@����?@�'p����$�q
1F,��U����|���y��1��+���'��ϷZ?7��}&S�bE���3���t��nZ�n��3>:��3W��o5$ݮ��7��M*��q9��^/�ϛ�Z蓙6@%#-�@c˴���z3B��<���<�g�����q?�@�&I���-`Xw���@�s�����;�
5�dTX8��{� ������S���뇌
�
5*�hL畬����O���:�ЎP,L'2o9i��!�t"}���:r�Η.!�;���)Y�{&�	˥�K�ښ�/��j9l�VP�mꜱe��`t/CN��l�v�X��J�ڥgp�G��V0�
��d?O�!p�Kw�1wo@b�L����L�1:<(6dtd��*kP��O����p�o�.ήb����S����`i�m�\^���9e���ch\� *�~�f<�͉]@��H ?@���?����wNM�>�J���噅���%�-O���|[δl�(o�YGa}�}��*��<F��������Mo��AOOJ	�FU��(�M���opaf�2��2�{�ۗ�-�[�v7��1���w�:�����ǆ14~�*ھ��߅��-A���ϠV���߬���N 54�D�(�����Iy�(��aɨ��
%�x3�Ux\��k�q�eEF���ˑ1�'�{*�"Z���8 C2����z�7#���O?��|��x��38|�:������7�'��I?�C�YۖJ��Q!��?X	��Jg��n�V}�=���[�|G�;��(�bscW�����8s��NFѷ�]��n᛭�m�َ*Z ciqN��gA~v�a�ǚ@Y�
n[Ef1/+&jX(�$p`�i�cǎ��b����������q��_VE���VB1�
%	�4�*���:�����_*!�ק��z����F���!� �������
j����2�x8�ɽ{1�gTS$��Z$5���K�����ƁSEd (P����c�5#�ѐѠߌ�wjH$"�.��tMU���h���_��~��Z�	�x�>����ξ�
{�ڂ6�J���c�NfH,������>s�J�w�����=ϻi{��m�j�(��q�V���UmS���rX]�u7������������g*��Fǆ�O}
#c#�˿�+|���܂Č =�>�11�Z[�S��6)��s�� *M��c�z�,�pFi���809�����f���Q�������Mn��(����h�(0f��_1�hB:$:��ȑ� �c(ڷI���u��n!	���A>�.Ϝ��l��`kkS�κ�2���7܊�/�_wBl� =�LOk��Zi����b�T8����I\'�g�F��j�a8xNx̤��)����NR9���j�ؖm� ^O�]����v��7���S?���ؽ\�	�g����籙���&�6��|�*��Z����`���k�̄�H�g&���5�_>,�Ơ1#_�s�zx}C��t�~�'�G�ۃ�'.��R�]���v��r���^���1�ãV�+8���0����@:�@;���pw8)���@��GLb���
��5K� Ʈp�f�����9�J:ޓ'O�;߈?����ӿ�
��N�|��	�kY��Gq����5��upt��2*���A|�;����<�"`�9?W��v`$�G������Fev�6���~yvq��۾��@��o[T���Z�����/�Q�S��`�#a����U?U42�jhammE'�7Z����Ĥ,�O����FP.�;Ї��g/]���<�<6�m\^,"5�S�O)��
�VC2�E, ��]ƅ�� ���zqK�H^���A�|\���zxI���yXa��UŤ��KE�k��6,P!x�F���Ȓ�'����ˢY�����8G���tˎ�����t�)M
����g���ϋR\�{`����7�I�su�%8򹑊�d��{1<0(n�l;X����2�;lrZ\m�x�_���/���;@����v�_U��M����j�U���۶r� ׶,Pav���M+����\�V%��y��(֤�ϫ6ӓ�D�1-^l���#E��O|
�Wm�8)���
?�F�6�euQl�݉N��e�̅�$��SO=��GӚ�⮻�҂����%T�dI$,vE玣�̕!+�"~�� ���C���p\n�Eg���&-�eR�����3��Q	]��Ĥ�m����%P��nN���Q��#�hc�54jTL�sU�)+c&��0{��:?#-��[a�����\0���y˴��T�VL��C��ڑU>Ύ��=��.�ͫ�	�5N����������}s�K�+ޠ�" ���j+E��N.q\ـgTL�NE@��i#�*�|��cCC��(�����@��v3[����aA7�X��@��T �_f�x�t؍�q��?-��a��Zo�]&L�SO"���ѐ���ғ��G������Zӱ�9Yl}��۟�Y�8a2�h��s������as3���."�ɪ�����x��k�QfECM�˦d�{��y	T(��u�c��𞵬�����{��5	d������6ڿ��>�s%�2;;��/}�~�4�܊&�G�[*m��Hi�>�L~J4���n�����F��F ���5�i_�$
E���L@��J��1��=h�b�+ͮZ�FV�2�,�JiQx�,��U�T�bi5*HF|苹q�'q��pw�Jџ�G��N���|&v�SH�҄�Q2��R-����2��Hʥ�u<��Y�.l�T�w�a?�FD�CȖ�2�#�ޗ��C	M1**�r�W��?� ��Tx��1��vh$��~����o:8�������?j�gv�0��x~efa��T�޸�J&���EJu�9�ܵ�]���.�}��� ���q��a�qۭr�c��ff���4�1u�(n��r�dr��4+i
�z����U���KX�5e�F+�?�L���T����.j�,L��f��Z9g�hx�F��(��o�C�c��.z;4w�
?�n�G ����Ye�۔�������U����EI66p�L�AoO�ǘ���/�x���͕p���������Ȥ������ׅh�յ[�ui_�ȨP�Bm3�^T�踙��
�\�:'��ҋ�Um��Fړ]��eK,��sE����T�&٘����eZv��woj��y�sT�?�����[���--���I��Gp�7[�Q��yYY�����!ٕ�N��prY��z�R������\�;m�zS�?�x$KVq��{&&du��e\e/Z߈ip3Fka��v�[����(ذ���ڙd��dR���H<lQT9��A�)�]�(�d@X��WZ���ylm�+{����������������9���GS�6�Ť T�5��X��2av����ςS��������a���Hˌ![�,ߋJ���Qlg<ٶ
x�II�J�hT��r��tn-¤�Y��y睲/`;��Wk��>G"�VV7-��T�m0���59-*�(W��F��p�i��H_�zR�/0�[m�mm�OY��`e+���Md
���$�fw $��h4!���N���O�t���75n�w�K%Q���3[r-��vx�_	7Kf��j���D��g���H�G٢�bӗg��3ψ�#�FƀY�~��l���gZ{��m�(_�l�s��w�c>������k��u�~�p�2�������Wn�,x��5N�>�3/�U+��K�"F�1t,��b�����}N��.�$�jt�km���K�s��q����j��Rz�dk��E�D 1�`z��!��N�r����O�y,6)�њ�.���˕�Cw��iM������
��?���%�ā=���A=8�b!�5�ܹ���K/�����W׭}�k���=��9<������1��A�]���<�\Y�5��*�Hb0ƍ��k7݄�ptm��d?,6�x�~�1�X��3�A$!��A�JR��TSΙ73�<���Z�쬔ڎ��eU��JU�7�=g��׷���Wn���;��կ���c(�9�*�x^��#��2S�`RܨV���|ػg~��[�㿊Q�D7{`*�ɏ����|���lV�����������	�F�@�+�´�~��P0�N����"N=�}��Yx:UD<�}���W��}�����U�2���d�:~Btեs��_��ll$�7���O$��&~��xc#x�9����7�����7���7��:��2V. ľs�-1�ZOmߧ����߈,I�)����i�^�D���"F�`�q�?%�1�׳��LF����;������ݽ���(�*���`�k��S'����
"�$�_}.-,cycSs������^��INve+�@%�p�LDcr����g���t:�o������c����r4 ���]^�*|�m�\�Co�n������X[)#[!m׶lߌ�������Fb��l��= m��ɾfg��طO�d;�Y�13-�>��c�����N@��57R����u4`5�y/̊pZ�A��{�6���I�\��4������,.�(苭$��L%8��J�V����{R��p�1?wo��k�x"��HFZ���#�m��*���	�	X�֘�17�B^�b�vd�*�
+�T&-͆��A2A|&x|r�fG ���V`�`���h�M�Πl�:4b��7K�s���A���v �yo���gs3ۂ��}�U��|>�`0��cq�M�17dU���*t�*����7d'MK� �AR�t���`�'tc�8#�0�l�x�Ha>�^���l�+(T�+���.�<�� W���O��c��#h�;XX^3�q�n��2�H��Q�&����l�b^S���t
��8{�9%�7�`^7��ԩܷWL��ʊ���J��_�z�~711���P(�Z[���~	�s����5a�_ؖ�W���8����c�(_���;��e�������b���s�X�����{��[��k¶�?�yf]�@�@�Ѣ94@ׄ��:o�=bk��x�b���l�3�a�2#c�ڍz�+���"����V���WB�C��64z�Tr��D�^���^��z���3c)�Ml.]V����$�NH��˿t;fw��������}_�[*U0=;���^cΗ�����`�¥*5 �qL�:�����S�,��G���!&�gװ�g�@�R)"����<�Y?�����D@�jgM��������b����ko�z�Ղ�RG@�^�b���>pO"�s��+��0h�B�A��=��#:�r۫���w� �ai�j��,�<���)�:w ������.�1s�z��V��v�^^n 0�k�Ą�,\��þl^�:TF��+�,}�r�S�� �vc�p�2_gЭ�h�jbTR�&�)!��C,�h&�����qۭ���;�����=���<������������M�,�[��eT����5-1E�DT@�^�h�n� '�^{��r�0sB����>r�<�W�/}E�
7���ݸ�����04��cA��C��ݾ]9��fD�kc7'��:\�B�^
<C8�G���<~�*���1*����ٟ��ע�e��p8��@���M�m�	�p���G#i�� �Q�=]��76��D%L��R�|/t�X��V!Ř� ��C��RE�Ό#=6���U�>��V�n�A�� >2*��#��)��	���R�DO�T�A�L:e��׊�,b��F��k�n��X�RD�Ss�<��o���V���k;})P���^?�g�6���MH6���\�u��׏E����f'E�a	�%Jo546�+
�6��l���ҩ�i�L�u��5-�mJ>�HjZy�dl��0!4��j����	L����$0#@��Ќ�ԛX/�Pjv�Ykbn-'F�� ��4eN*���[^�V��
Eb�i�n���dF��u�9:���9�UZEZ&���N?�,*Ւr=,���^t�|�
xRC��1����;q�����5��9�Kvl��'g����h�{^/�O"�Ӻ�z��-ȴ`¶�Rs�-V��u���	���tt_�},�J,[��ku[J�!�bl2-jC��r��P��.Jȴ`�1"R2+2)��j����|�!���5C�L�Xv�ϻv��Ď=��HMD�F?0��'�r{��@P,+�t�b[VEc�.�"A�;uԪ���0vd(q��x݈G���(��a��32��������&:�������SOJ���3���%���v_z��zk<��.��!��z�9p-�}��>Z]�V$��l�T2�Dԃ�o�:\鐭�Q	���
�~x��N��t�������e���窇7�{��m��뉻T�� r�6�_ZP��a�A�����N?�#47���U��T��vNbj��Pg��7�Ź˲���C)��3i��IQo��x��8�/�����O|V��nx����Pi2�:��Y�b����Ȯ,b�o�G�enśD�f�G}kιi��c�B_�dT�Q�6J��;5T�5�~�t���uU��q�H3fpL=�;��U��a*��UAI��׬�h�10:6�J�����э�ԅ!��ߨ�):z1�����@��S�Y�B�L$���ܭ�8�!{�=�s���
�����'O�/@��=4D�:�vñ�+��7Ո�Hl5�u����u�LQ���vpb7R�20� ���`:�o,P������>g���#���
�,���VVL�kNטSy3����	�����֚x�oR,�SO=�P�[}�S�0@{1�f���s-�*b(x;n���8&wNkp�1���" �L�9 8D��9:��-�L`ia�	
k�����a����MQ���J(66dn������ ���{l�WLɴ�`�"xI�g���\��s�y��Z��z�|��LKO��a�z} ���?{��֨�½A�FE�%��9 �&�4��yi%�G��PCsX���� ��.͊ۅ�ߍ=c�1��x<��ф2�؎�W�&f�D����f	�jSA���&���1$F��l���r��7H��,�\�+)H]�m��H7`�l���"l��m�*F3I��$�0˶�p9-�K���/�_^o����<��ko�a6�V5��]Ѩ�ܱ�z}��Y�m{�yMg�6�riC�JL�cQ�ϰ�>��ˡ�g����!�^�'����]iۃ����� a7�^F�s��Ɍk���K����7\�v�a!�Ip��U���8~'���~(�F��}�Qq�R�=xʭrUZ������ߌ    IDAT�%@%b���\C��a+�E�O��Z�$6��M8^�n��Y;d��ha��̝=�t8~hJ����B�h7Z��q\Zg�r�uR9�������q��W 5���&j�A:��D�F2q$��2�5�v�ܬz��p؃{f���F��nHd(	TM�����w�'_@��f�`������Y2*��?�FǏ�b.��Q�a�a@�WΚ�ݩ��ٓX�x
��
R�<+�7�(�Vߍp2�D&-:���F	�jU%4N����e.�����"��O�-6����j�~n_�D�kp]GV�N��A�Z>�R���:Ԃ�1(�/.�����p�O�UP���z��;҇�#��[үP�
�9e��D]S���ß���2��J�*�#�HgF�Y��9p�r�2�]�������q�0l��X� g)�Ũ��z�q��K�BFE@��3ŭy7����B���˶Y� {�`�bK����}�(��P�n"v��\�k��ǟ��ܡ�-�j6�YqH�њ�.��5: �7�k�>!Fef��Vz�G������k1�.�r��a�ӡ�ԫ*G�K	k��D���Ϫ�'mS?����Em��I����4��k_��*S�Du�uxc1�����"��gST� 2I�t���g�e��B��Ro���B�C����u�Y���m�*##)��q�\VC/�~��1��_"AVB��W�X
p<x*�Ri�]h�=ddth8 Ǌ#�hq�A��v��4>+r�T08�+�Ӷ�u�ۀ��A�j��EB<l#*���u��N��+!j�vn�!p��H��=��4	��<p;Z����l#�9�@����q�3�i�DCH���;���X�vU�) jLJ�>ί�c!W�f��R���ЍJ߅��Y�RA3;��T��S�J� �i8b@���O	ˌ���[J�����od��(��_D��M��=Bul�0�@E���+��5��^��F����#�7�Y�I3���r�X0��i��v�I(�ң�{��e��|o\�ml�g/m!�"Ų,��4`5�;h��ט}��dV��ԱА9��j��++7�of%˴�1	�8�"�r@��F�����H�䑸���OLaj�>��Ď�נяc�쒘�����1�.Z﹗����̓��l12X���'���ֱ���F�����0;C=���A�J���h6Jz=�M�O[6���p(*=F)�@0�ə}�u���4��(�u��BΨ��3�˅d܏L�i���Zr#u]4�U�}����7@�{�#���v$>�Gx�����Ri,ֆ<s9�֎;&F����b�//�Q�]u6$.� �C���Ο~�g�ZA��@�����xH�s&���V`[�֊v����{�^8z�N\��7����ᅅ<�M7Z� |��*g���]��k�2�k+F�D{Z��U��89���>�����4=���bШ�V4�d����SQ[K�F���n��f!r��z�J�$#D$��d�c�tn�t:�Of�ˉ�M��
�:�2��
�QƘ�}��Ӄl
-o�pP��͍��U�a�u��MP���*���J��27@>W�������=���j� ;Ӗ�W��<|��w�[��}���B64���=�"j(�X��d+&kUe�7/�H������J�3n�̧� P�#������q�g�J=��2��V��T�089�S���77%��q��#1��<�)�ۢ��-�ddF�Fq����q,C�0�n�e��=16�����#e`��%慟�g��`4�s/\£��>�Ũ���%��mJ7�s����� 4�쪥2'{����:H�X�lжz��`�*�)7[v��-�����8�qQ����:�k`iy{����h���\�Ȝ��|}���l��-F+���۟G��?�pmPo�5W���Q#b�$��E�B��a��"�)+�QN
(𳋹q�&��@�Ɩ
?{��F����L�Hɐ�wM��ɑ__�g�(�[���T�a5W�[�:�ΰ}oSS�HgF�sv�7�>wZ,R����Xv��fz�]��FB~�٩mueI�5#�9P��m��m+MU���_��$���d�xM��ʅ�t0���������#٢6��+�zV�0u$�w	ha����q�{�	�|>�V�µ���aЬ%ݲ1v�v2���`�(��vd�%8��&���	̶���|�����0��Ř��4fFEl�F����̮2k�/`˵F��������F�3�� w`�:sz�`J�O:���</XpQ��k7��ڥ�qL�&�B�M�%wg���hԇtă��Ed�.����$�o������I 恐'�cq�Q�N�`����Pk ���Ge]g�"VLL�-F��4�W�oړ��H`�ۃ|M��b^���Y?0����~�=�xYؓϯV�:�����o���o�r�6Ξ�G�������'�t{L}l�XX���3X�{���k#H7�=N��mؠ\Nd���[��b�v�����,�w�A��Cs@o�a ���ꍶ��;�h� ��!]	�+\��)l�29�T7�����p�먗7�,��Yʣ�*�=�h��k�hٖ��x$�ʟ���3���ݘ���jH��"	G��L�%��ݵ)��P}�tR> CMNv��Hs`Zȫq����� �G��1�!Iw��~��x8��.^r��m��9<��Cx��9��!��R{��d�A�*�f���ي�V�L���ҦF�eA	U�-CM�Rb�se{�܀u��R�ӒI`B������������{?����z��CP�a�1�@�~��nT��ҟ�OG	��<�	����ut�0�#��@�PR����Vt֒����i��X{���ޙ<��7e$����o��Z]���obeuC��1�Ԧ����+*6����R�4�/6�W$2e/�q?�<\����3��� ܋T:����E�1�=pP�CfEbf�#-����1��e�Av�j֏�0]��D���*����ka�\�붃_>o���̛9����r��b.��ϵ�h���֑���~��P����j�-\
�5�@v� 66sb�����Ϻ4*l'�+j�Pp��֐�1��a��(���xa:[�V˵fk�
�7�X�( �Y�F���'�
YZ�S�;�w�!Tj�>󼱑:-	ZA��.1�^�L�_w�<��s8��ILL�)������)�nj�bk�@�2X*\C�t�x��7��_�:J�
*�2b��Z?�f�kY�g/�+i>L�P��6�9^���>#v_�m�)!0a�����	����e`A�:�׈܃b�Mۑ����2��O�-5�7;L�6����a��א���3q�[-AF����֏
(�3�8�(�o%����aK�b�.gǎ���ދBh��&L̠�I��.���]�BS�bX��f
�5J��6�28_�-`e�p��Ĕ��S��#&?�"$SGas�n�뫚գvL9,R+y||J#Zb����6亂�}��{j��\Z�������� ]r٫K�5d�!��3�o>��XX]D��Ð:&>���N�Q������:�k~���?��\�@���:Μ�S�=���2��E�SM�Z�b~/<��::�t �p�	γa�$�~� 9��tCx��gF��Bzd��BI��6{n��5Dʪ���6)�\`dm6���lPUݗV��%R�\H��8\IO'1;s�n%$P���(m`Ь���,���Txpr�q��#h1��y�;*v#L3�oF&��
��o�t��)"�͕�k��M���lr��`+N�����W�XeuMo���ɂ���Ll�뮻Z��1`k��jj���C+cÈ$����-��l;P���hԌC�}b������N��?�o��AP����XN���l�CH�B��@�v\jT8?����/��O~R�.E��HL)��d�4=��(�&���m��_�c��{`k��.+;�����hTFc1�kr���*W�G�9�G�R�?��Ͼ��8t`?��w�IW�����[��+�$�x�G?�������q�j!��"�ˋﻅV��Hħi���t�H;
�}jM%�)^O��t���j2Յ]{��g'��v�j��d��U�����Dmo�Y�>�9A[F�b[:�U�U:5Uv�l0�<i�Ae~c���������!߃	O�7-��0�>�>3�Ť�D��jנY���"$c����@���d���]S�MF5ɚ�[��*Uۨ��J�^�,�Փ-UP�P<P$�R����=SٍM���q?�RÞ)r0�i��o���<�y�$� c��F	�5�_�jE�������s>Od��|�o���#��G>����Z���p�صҌ,����;�wCV������ؽ`{�e����%f���G�����𗲈�16k����:�{�H�׊�
ev}�3l��I� @l��~�'�fK� UZ���u�?h��\aS����aY�=l�Rr;4��;vbv�a4�~���c�fU��4Zn�lro��q��NW�-'�s�T��6M[��|�d
�������p�X��d:Q�1.�4���|�� u�q�odN��zCJ�PqL;	C� `6t��X�楅#>D���H�� �J#� ��݁����_Y���BZJ<������_������˂QYXo��5zx~n������4Z=��=7��i�.�>��kI����4��-]l�-ce�6V��+�aN���7�+䟽p�c��Hm��c����(�r�C(�D���<�9"(�(����Ȳ�(�=`e��*�5i�@��p��J5��zq���9D���C���);�N�΂U(�)M~�A�Adpv�-m�A���ai�-�Q!��%P�M"�R�cqi^Q�r�P�(�؍H(�ݻw��[o��E�os3���E�5��p���Vk6�D�xZ�b7"����U�$���בQ�+`��f{�|=��ww����lٞ�u`�pF�c�i-%̡w�{n��=��@�tZ�'�}�5uz��
"�"�%]@C���WMp�㳟�����2d����ظ>ת3;g~afJ�9"��ͤK�R	����,�[n�ǯ:��<�0�{�� �������Xj?��Sx��Ym{Ͷ�ذ�A8藋lzbL�`nc� ]!�k*����%4==�;~�Ny��q��9�����qۜ�<:>!����<(�>�ƶ���C�F�T����e��&�^Y��v�վ�|,��W%� K����u ���ܙ�P�(ʕ"B����o̼▛5��ԩ�x�[�B�lrZ�.���*@�Qa4:5��C���qô~�~*��n���b�g'�09�D*@��8��z��j��r��|������%TZ=�=t�^9��<�S#jMq:��O���㑡}��kp�"�}�oP�w�6.]��L*�����/ ��*�'W01��73��[i��*��׾Z�s�
���ra��CzF��1#3�ަ�*�Uo�����m�����U��=�>Nk���찂֜$cˠ�ٯ@s���U�L��R����E(`��v��x��g�wq/�@َ]0,�?Tx�p5��բ�X�:�s���{�qS�ybj{�A��B��+2�pf7���}�P���V��ۦ��kȌ�ЬVШ1�Ss�p�g;�������jY��ѐI��4H%9P�g@��$��\m���\��3�}�A��W ��C$l�C$xoy���P�tѬ����4���/��Ҝܵ��\24�{f���x߽/�2_j�.Tw��[���0�q��6�m�;OB�&u�J �o�=������Ѩ�Pέ!�]D5��f���2	[�K�)��#ȌOjS�Bz�(ר"&P�a`�,a<��I�JY� h}m�zA3���~xHq�zP4 �1@�d�è�
�bT8'(��i��a��� 5�f���Aea=�z�f���M����l2���'L+�:�X0ׅ`ť�z-��cbMJ�<��/
(�`P�{⦣�wڨS)�>}�.�O��؄6.n҆�7hH[Z��4�*���c��{��F{���_k����՞s�����֏= �symY	��4@�lr T������3��3�H,��ך�OLK&��dhg֏*ZkN��\qS��g� 4�3Z�͐�x���O>uRɘ*r@�y��Aae�J�sS�"v�n�y�fҸt�T��#2:1!m�S��å�y%�6�5�f9�����t7_-J�M�|��pn�ʚ�;�j9�v��)���n�፷K���xiAY'O>��=�j��P!����꺮�˵���gF�^�n�*�$uM���n���B!���'�m���������?V�< m^�e:�eK�����i{��	�]صk���������򗿦Q�.-����-�g�.��#t���q��u,P!s���^�W�1��c��)�L����c������z��\����"Vs%Tm�8�'G�?�0�X"!qc�X#G����������>d3N;�׿��-?�^8�QLN���3�N9'�8���5���y�k��^݇j���{��E�Q[���q��B�6���C��'�r4H
�9F��7s�l��ʟ���,дk�@��0A�^k�p��]d�N�{Yp�1t8��-1;����Z=��(���Hg�׾�5}N��p��.��@Ŋi��1��̻!�Y�n��41��s�d}(N���Y;l���V6r�0�-:�-���9�U�fo�v{~na"16�A���Nð��A���uݽ�ɱ��z}��$c11��[�b=���X��T�q##����>�� ���}=��*���&�j���fޗ���aG���I�}ؿo
<�U�-�	�q� 1���{��������F���������� Ŵݡk��_\@��D�B�q\7�lbԚpZ'�G�-#�A/����V��54*E	�\�]n��hD������j��K348���;�^34�A�*q�|��	T�+��JbB�L��P6�6F���������)B�]�D�V���5̰��h��P��M�H��g�ٴ�T"6��T���>��ޕF]��B�(��Q�;c�	Tx`1썳�HK'9��ܜ���:p�͕�az�VWb�+|H%3��Z��7i�`q�9����l�k?�l�N�->~�����>�V`+1YS���|�xX�f�h{�`���*&✇��.��F#!��20�.�P�*�iWTO��g��p5~DZ)�5�4s?^����{��%DfFEǬ���R��4Pw{�����pc7 ��~Z}���
Y�:�U����	�8�O�z�X¥�y%$�.W�k�[��]Lf2���~��e<���J*\(7����5��u�|Ǯ>����wp���h��b	/������8y�
�2��Q���]3,�䁹�<$�Y�3K�cA7�����z�5���7Lm¶M`(p�d̿Sh۞��bF$���C�T� r;�x&?�ݨ������?���cx����~��^��n��oOH�D!*+Js�:����QRT�`}$���-6%)zH�I�'�f��Q�V���O��26,�"�̈͋�h6�X]۔�z�F!r�)�U��W;�#�ˋ�ޣ����02�V����r����5]3�B_}�m���;q��7RaL^�'���o|���/_��奬���eS�hڷӦ�=��R�i�d�`�ΆZ'��7���z��u�@�-бe��I���o|�	lh�U;�A����U*##c*��:���?��	ԏq�]��E�Sj�;WZ?���1@�@�ѨXFŊi��,pf���ʘ2N�y���zUӓ}�݈�w��K��v�O `�
[0�|�A_a��d����'�Ѯbue����m���![�ܭ�����|TT+��c U0�l��Z�gK���s��JV��!�o�R�)�|�0vL� ���˕����t�N�jA@���]x࡯bn���:O�� �~3;�#v�?�[�x���������L'��*weK�0g�0ve�����P�vQ��	0��6^��6ï�!dUe�7^êZRS-��ж���!    IDAT��Tmd=��hu�]�6�_�Æ-��m�5[t"�����Ш�Ą��Pq05I���R�L��p�NC�/{�͢f�m#�u��IL��5I��>�Y���C��g���]�e�^�]ir(3z�@	��y�S�ٖ���L<�~%g#-.\����{&n��u!�
����pD��z��ރ�ꡧ�D"Vl���f�T���7�yO dn\<��u��g���K�������l�}�| m%n��X�^(P�J��v��DVCw���UL��k�lw�&ۧ�7�T�"�M��2?Ԛ�H3S��M�'�P.?#��[��V�3�z��_�s�aq��x���X ���f/ �qK�*�T������cjf*զ��y�H"ѥp��t8�;~��H���c���HL
s��<8z� �{椀��'��wމ_��_$�}���b~�{��|k���I�o��P��g����d�N,�d��ַ
��b�=�T�g>��s`��� 0M�u ����ɴ5��t�H�J�G$��F���H�C?���x��%�L&8%  �V�a`�y���~^
T0h+Pqzj�� F���d�ϧ���j?jt��4�XY�cy=��j��	�|XD�\��: �?��#s!-�n�{��W�?`mm�~�;X]^F"A"�Zv3�f4�L�S2~Ǐ^%�r�+oְU2�\����~�Q1��<��k9�K�Xjڼ����;�j���ٲ���.��e[l�PNd���-c"4�&ߛ܃c�K���ǖ��*t�����4�"�LxRgw������CL��	�3�=󝶞Ð^**���1�)�DL�a��7~/[I�^a�w����#�`9�Ь��/bCJC	�=�G웑�/*���h�x�r�Z!O�z	��x�ր.Ӯ�Nr�V,\�+��+�#�`�k��9�|fh< uE�!ǃ�{8.��Y�G�w�a�x�^�hi�E���a�ci a�9��ݥOT���v#� �:�}�~�p�<ZV.}i{e�L��䃿��k�O��OO^n��}���b�=k�N���G�2�����f���/jS�"G�I��>$s4�\4Q��~�=����6ՖA�M� ZW��9��_#R�2`�LC���M � �6�7VШ��Oa����?T�#q��O��~ 4@˿��~��n� ��ѠG�A)�gC�>{> j�Hlk�Z�\�.^��
Em��%T���C>VWT�^�Ne*�����Ш��bN�k=��Pn漖D��&,봇}��SF����}t`Qhh[?jal��j7+��b?3-�Ač����-��bg�c�苓��&j]��MOT�s���|pN�����V���;}�T"��xz�׬
=^�Ri�(��":�
���bJ$�j�8�hۓ�����Ú@�Ο�����
jY���+�gieO=���/���j�
!��Ё��N��9�H���/u\���&ds,-���h��0�~�rD}Z�����M%���� ��8u�)��-9v�y�o�u��CcP�,`ii���c8w�<V	T���Q(�k�uG�Jk���k��3s���f���W�7�b.t^2ٶ��@,Ϝ���&%S��]Pt5�EL���ԩ���g��>�a�OMၯ?�����~�����#�1\��KY
�:|?߶�g�����O���H*��SЖ�1=1"�J��"��![͕f�Z�r�
6�,�����ݔl����G,x�=ABt4 �e2��S{�M�#3��3'���gNcb$��wvE�q�\ɮ��>���x��ކW��jK�k�� �+
`��D�����V%�����0DT*���#� ӿ9�2���=�3�R�])N�9�k�,���X�}�ȏ+C���{�G$R��~�+o��V��=�>��O�_�*�����֦˫�ג*bM�Ĵ���\�n9t��Ӣ���5jCk��iHd����ž�Wa�Є?��^��$ܡ���tMѽë
�#��I��7����UZ�@,�vi���ׁn��~�p��r�#`qLr�If�5�)|Fy�� �B����3�-�kc��&���Uhu���8z�qBL�!O.�r�pqDE��d�-F塇������F.��F�viqf"��?�����_�
�J���<�V���B;��Eus�׋XX�*�-�͛����l�5�l�(0ٶ�~�VR�k	\�Q��������]�+i�"�j<�FbnxÈ�	T66�h�*��c�M�ƨh�n6S.����J�QB���VuS@���t*�񡢠I�C����[%��z�Dų�#��V��k�T�5�4:mmd��kt{���u�����x:�� �Pa��� 8��|�2�k=$�&����cj��j6��5�[m(;X��.m��e5���X��ZF|i�S��~�� ������I?�z���0� �щUq�)m���g[E|}V�:H��Y �ƻ�Т��k��zK-���:���Vu�(P���]�4��2�'�jN�3$��i�O>���@ԿhCtz��XDZ�D$�kN�xfDI¬T���_ɑ$���V'�=���5MB��ZW=���~�7J����E$�Ů�)d�� ��ɟ�D����x���o��x����ay~Iiȏ=�],-�ay9�^w�C�0>':���S�2'mt9[1���zv���ع0��p��`��=�lu��4����yrt��Y�!�V�ύd�n��rT������C1(_������϶k���U�J��ɬQ<I���*+!��PQ��Îi֩���fv��N��ov&FR��5�G��B�T���l���|	�z�VOs�FǦtH���8�، ��~�f��B��0NIq��^Mz^�|	A���N-Qf$�R��1#d�|�P�_��_��7�R{�NG2iŊ\}d�9q�G?|R�bz9lz�`d!���g�󓢑����*ֹ���W+e[؟/; �%�ϩ��T�\�����T�$k�/��f��[�Z�̇����g>��|�+���&����R+��Pl�8�o/*�H$�Ki�D��`�V��6��ME��Y?с(�w���F��,����q��tx\L6�]j�LKs�
E��P�dD����<�&���e�WzE�i�p�D�)*�幨H|V�L*���rj���7ɨtL�AJ����'�1�A�&�L
�">2�c�O(��5
���B0������.�F�I���x� �i����˗������?�� *��~��Ͻ�tg���Fw�� ��6νp�Jg�;�s��C4��p@j�T����!Tk�r�K0k�%��V�j��M��KBU'���"K
��������������6skhq�e�;A��IT(�g)�LϘB"]?�4JY�8u�[�k���._Μ?�>�V0��jkU�]� S�υ#��4٧��T�ː�a��L���ؼ&R��(v=FF�=���	�h]��iD�mz�]f�Z�^�K�����D�P�_�|�8~�(d�y�E��x�,����E�bc��0�߶�,��@�Ve6I� ������ic����Z���@��$�]Jy'o��:5�&SB-6�G�\�e���GO(`�O�ԁ��'�zk��Z&��٠hh�#�4/I
�A���ЙL�VX��`$b��^�B\�dP����Wd:�]}���ju�����JV�hSm���lAF�>��5���kK�F}�+�Y����4y�
�:x�0~��w�7��>a6ƥc�����	�$P�v���Y���s�_K�I-?�̖���%w(�VX̨Q����k�I�FY`�u"������X����M�_�RY�?#��FVT�e����������6~��~��ؽo��J�avPH�/��8�2_��a0bH���=暄���=��c��H �f���,��]�m�ya���h��	��<W�XY�@��|1"1�q]�&����Q�ܕ$T4��S��	��H�(���A.�!�Y�B��8�c�N���rzI�`<�o�%����.�5�����\~+��Z�
���[<�-���H��ͅg��]'��7��ӒQ��<�������K�L\6ϕ#.v�A&��kN\�뮻NQ�tF����/�o��o���bڲ���%Y5e���cD�Ԩ���F�'Mr1�4#&�X�������c�?p_���p�ĺ@g��F������1��+�Vϧ��QŻ94Q,���wuF3q�ԋ�����ɷZ%�_�H�?��u�	������Ϥu>/�?;C�G2����^FE �A��C&��F8A,�Ğ���&1��4��s�h����Ѭ"ra�T#ct:vQ`�n8/r�������������P��ڜ�����̙��j�Pr
��r.��㹧����X�nU��az�T]�1j������֘m-�>�o�h�1:n�&
�C�/#�2U����#Wct�E�1��5N�BF�:q�Z�PaeL`@F�㦷�C	7@�O�@�SӼ�Ŵr�h`���9 %"�J͸�L�ߛ&�R����g���X�BF� lK-�$��a`�l�
��VW��"-L��P,�*��ϪtrrB1n��&i��O
13W�̊ĉ��{ p*a�$�b��[�b6�1� �d,������lג���)�~7��"2�� �-=ð�ÂY�DI'��¥���G�cv�^�O���Ϝ��򊱻Sg@q�>� n��T\�F�d<:]�7!���$�{���觌�h�����66���qh^�#&��6�+���G��fW_w�2�hm����Ab�GզE�X����i��TLbZ��dRq������6�u7\�����ě�C���u/\���/�ԩgt���-m2*v�m�:0��R)[5�]�(Ez_�#��}VeKk$���ƿ��@V��xXn��1�e�[OL��/�O,�0����_'KH�2�s'���cx��އ��_��]�*<���k.�֋B��e��c;�i�.��.x-D�.$�a��8�A�wc��4���XL��鬠Ey%[���
W�����F��_�us̰�I�2�U�7�`Z�N%,D�_OL?g:�P2m�����i1����)~X�197��u�\/�
E�zf|G�G��'�|�JgN��ٳ/1��aB��R{��z�_g���,P���M���~�e`4V����O,k�M�9��β7���u�>R�|�kN\-VsddTC�\�}�ݧ�km}�x�a����@� Lm�-�b�[~.Z������1��s~>����a��5K�=ֹ��#X-���L�:L���u���3*��#Z�M��-�2�!�� �NI�J7#��.�}^w=�Q�^�� �{�d@l�4�s��x��c4Cf���>7����u�(��E���} 3��4V#K��#�� �����6�*�:RAfv� e�ϕ�NB@v�Յ.-_<��;��[��'6��7����w_���g׊�Z��o>u�򻆾���`��#�o��y�KU<�ēX����UX� SY]z��f����c�$�Aߍ!�w.?�Եx��2�~[����b�����&�lV���zh\���t�8
i~/\����	0�l��Wx�?Z���V\P�뇳>Ȩ�]]x8��⼡�6�L1'ᄄ_v3��n��`�]�54u��"Z�~Dy�v�Y�������L8$w�iʉ@�JvmYm*�D���-��L��L�O��?��o�b�b|��sx��b����ciqY^#���uP�j{�m�b1`�TTv��^a�V���m��2(�d�5Ш��"P�'+���Q9Ȏ?�;wb���8z�Uj!}�ӟ���E�B�h� 9�ɩ���������/*v+ׁ�Tۂ�U�V�D�1�E<���N�zKKK&H�ܰ{�Q���Rj�2�3I��o�����������c�����ނ��i|�G�����S�g�*]&�D��>�S�+''�Z+j�i����I�
+�w��=���o7�ۅ�g���>}F���z^� �}�3P�6�কW�2d���)����P�mC��ѳ�4����fc�j��%��;�ae@�)N�o$�8СLa2[#�jE�"�g������@��>yJ,�D� �l�nJ6Cn#�#|����?K���I�����JI�1=9*��ό�RL[*�@�Qdʢ�����:�se�Z`���3̙7�Td�:�p\�H2
F�����Q���E�H�b*��kf��e���]�Ϥ��1���w���b��M�oT�x��G�mwT8�-�yǞL�$���d�N��9�'�9���Z!,�޲�����;v=l�5�)st9��V�@�
�p�	 ��u��!\{�5joqO�S,����^�
Ao0l򜴆�ŖɅQZ�V���O�҈%*\�*z�d�i�gণ�"�Ȩ���^���HOb%ߔӇb�@r}/�As��]�"�k�גBV�%�w�0�I��hU�:Sa굢��V��M��򗏚����x��dh����'���Z�7B	J�Y��c`$�{Fhm���x�{ab	:�2���2�-xe�%�n�f��F���&�[�VE9��8�o|�����{O����Tί����x���ν�� �R���z]sj���;y
��/i��VZ--���X^� �^n��v�4��iZ��!;#��x���!rN�[@��?p��LL��l���Ȯ���8vA�5c-�J��
�^��Qd���:��Td+���ߡz�̆!����z:CF2N���C��i��|�(���(��z�\��|<�-P1.�
�� >�@@�7��������V���7ڲ�CD�<��C�w~�=���[5J�����a],T��݇sg_���s{x�3(L�߹a6�\�+��`dC�;)�ۆ�Y@��y�$^[���m+@"N��J�b����ȑCz�WS�ΝӲ���C�����j��/�W�zҙ1<�͇d)�jgˮhrT,=jʅ.|���(�c�m3����n��t Pa��'�4R���sZq ���1���܆���7��^�s����s��^�ڟ�M�܂�.\�S8�xXpj6ZģQ%�9����g�*���.�����5�\�w����_�es_�^�z�I����ҦL���t��\�UM�{�^s`����Y:�j$�f��Cϫ�s�������������|=���?� ƀ�&1m`28̌H�����'�~�~��:�o?�]|�C�OzJ�_������?�@�EX@e������s:������@�D:��3�����hR��q�!�d�B���f����Xެb#W�>�k�C���XAz4��iB�^��qs�3xz�(
L�����eQ�p�nW�m�+���9���_�s*z���*����Q��	T�,1�G�zP�� �9��p�k��N�gL���=���C~m��mF�;�wz�5���CՈ��^k��5â�qtIm*ԉ1R�{�����}XY]Q��-t��S$N�b�ہ���l�{�h��Ad�C
Ǐ�E:k�ϙe�Ud]���$�g`��F���0���nY�����w9S�uS��B|M2f*�l7ʚ�L����P/jU��H��i���G,����dZ�Gy^�ҙ�5� X�s(a��R���L��L�����Ӽ��y� 1�D��T��,:�(Z�z����V*{"���TϞ�	�V��bQ�v���:�	}��}�'ny9 ��k�]́���詳�&��}wX���.\X@�P���<r�5��v�H���e&hƸ��1��4/'5������	N���a+�>TA�p���34�V@������AF�\����(o�V�e0d8vFz{�}2*��:z��P!6DO"?��(���5	ctd>oD������O�4>@���eC�с"^�����Lؒ�Y�yE-���@�}���4
��w��ӓ�-�(d�m�p@t�=�܍�n�^h�� ._��U�+_��z��\A��e9�PB@�3)��c�+=j{���    IDAT�m�e�ο��f�N(8=sU����~������}�N�]w&vLar�$F'���?�я��ۀ
��+�X������b����n��;"m�� �LQ"�������D����sЈj�a��֏&@7[x�+o���ſ��x�ϾVX���e����ƛ��#���SϢ���z[�=ɿn�,�(�J8�U2j:׬�J���଺83����]������oy�*��x����> v���D�t�5]5$��a7��ZN.�/1Im�uo�+bY���5�<H+�7t�T��q��G��ҴeG'A�dG��iɨ��5�N'����7�|3�����{��ӧ���Ϣ#�m���@���
"x�x����JЭ��B"��̎1�NO"aj4�����S:Y�P���P�N��lJX�59W��F���#`��K��si|�ԙ>���,WR�6=]��?�Zbj�|�A���f0�тq�mG�;�����G�م�"��<p���iϝ��˸~,Pc���"�>��Yu
��z4���~�2��Y��
�@�v����Z`�B�E�Q�h�9l�;��9*|��������ݥ5�b�3��k��kC��x�rs\e��f"�؊��9�X�S�����i���C2ώYbvv7v8�Bm�|�Ol����J�o�g3�|.���;����ivS�\�f�@�E-��-=������hc�k��oɅ�e� P�gu�2ٖ
��+����G��:jx �_��ې.l�!���ӗ��Qa�{,�C"�^����A�FQ�;��x�'���KP� �XȽ�o:���/n�7�Ϩ��=����s�&�|]�	���up�������xQwM`e�%�Ң�6b':�����ZgH >!�r�Q���^	i9�FK�AǏ�&g�8���fz��P���_�9Ș���[/aT��=�rFEs~��h�r[�D����3����)�����fM>����<��f�7d/�V��k����S�m��V�z�Os[樤ba�Ky-R� ���T���TT�]w݉o�Q�^ݖ�T�\�8����'���ŭ]gz�m�lہ�ӂ~�F�d�X:ײ%vC�,�*��E�V�k���Xi�'D��I�uݷo�t8;&1>�Hx�������߉��˂ 8��ξ���F� ���
P���*~8m�,�K�0	T�����l� 'ղ��j%��9��4=Ŵ\��r7\s�y����3O��o֘��.��;�,��c���˲[��}i!X�0����c���g9�(W
ȭ���B8d��Q��_��x�k^+ ���q�^�!�e��U��ݾK�l��g������rV������|}{���}��'���&�L�e��b���bb˒��jж���
7�%5*|O���'�����Vi�������Ҫ��9P�RN��D���  ~N��$(g ����|��î��H�"r�1W�N��Xt���Q��,����r�(ϯPb�"5w��>�A0���M�$�0����6�l�Rc�J�̢�|c�M%�8|���]x�oo�W~>�%�~�V���dN�*�89�����%@��<�֌`A$�?�ג�L�z46�L8E�3߇M-��kuLbb��,˴u� ��/�����d�����5���@l��zV3�|>����@XG��� �R--"\,�1�{�u��~8	�0@�0ƙ�q�?t�����Čf�0B��5�[��lr��hKq7�O�Rˮ^��Y���$�3�Q����>ztz��1hUPɯ��(�g���{�/�=Zl��cFo����#����n��A0�B~�8ݛL��!C�i�;���D��B<���	���ʈx���H�'O~�/�+��G=�������O�����������Q9�m�n������"�B��8��B/�p�fG.U�@NU(/�zd�,��!A^OW�f��f�eƠS�A?m�/�0j5�1�#+ �Dz�j0�ݳ�� N״}F
�h髕KҖP�|��CŴia���<���R+����j�65*�rZFL���L��#�J"�!W���#e��V��M��h�0��h������E�R�W��/*ܠ;uEz'"&�6��!�N�ll��@Q�I���]�z^��W�MN[����kXY^×���xꩧ5���X����{pZ:�����0�`=�/�(����߷ov�}�ݺ* �9y0�~u����C��g�.U�̮Y�M�kJ-��>t��_Ժ`vJ�B������M�3ke�3�'6,�f�p�3aJ3E{o��ax}D�q}���&�V����p�V��a�0C�J��U
E���/�W?b��nS���5|�;�IL�ds3�ۏV�,ǎ��@�c(���"!�_��6@8����/�b��2R�tv١��ȷ�rOp�,.V��\:8���v�g+����]4�um �*FWp%����F:8�N-�&���a
�D��h�m���B��j���=}���S����	n9N��ð�#E�w�SY�0��a߼M_�jF��1�cc��Z�A��WK2U����R��R�!����R��	�Ҹ�#KG{��/&E�m!�6D.����pH����F���hPq���+f�h$"�Կ��_��^�:�KJ��t�2.^���yK�G���-�֋3��LMf��3���V��XX�ӎ���^ol:z�V���3��c��N�5�Ľ��=�o���c��mɕ��i���ț�s�sh!��4\^wè����h�s��!�Ȩ��s�/����L���	�f�_'=2�=���P�R�/��O�A�j]�~gjc%;�������F�.�&����cӒ}��RWW��艀[N�fi��;��ځ_��v<��W���Y&����ɍ6I��Q$Gw"5��Y�3�X�pL#2|h3e���^W�t��\=$cl)�2t���z!��I�������#�$��@��we���~�_�,��3���a7�O<w�]�Դ��	�6��>s^��<jc�����u 0�w�Se8���4� �)�ˈǒFPD���%�g25�j����M���ՙ#aU��T�c*��_m�$�V
Zt���0�l\J�uh16�nZ�kr�����9��ѯq�W��dZ:OR�,қ�Ev�ܶ��A�vaffF��zS��ׇ�(̳@��x��&�m�Qq�J*�F%���N��j�vE:8(����q�7�|��]�����py�Q1����>/�RR��yK�e���kM��2��<�fc����|[X�_ڿ��=�,�bA����6nn��/(���q��A�T�
1L�豣�N锾��?�a|���?�2�<tZ��5�-�#	%��騴P�tJ��|��-6Ȩ������Y�3ܸ����}b��L+���P�0j��R�
7�%옘�޽�119_���;x���^��R2-�K>|-2IdR8��
��Rq,ˮ.)��.o2�܉㡘X���$b^c>m��Äb�\��%��gWu�e(�qO��֊]%�v�Y�t�0 ���ܤɄ���e~�Q� Rp� R�N�XD;����(��j/ ��T����(�vO� +�4M2��1��m��]�s8Ԕ^�/-�a_����8�F���;�γ�ާ�2���b[��16�6ŀi!����	\ @I.a]��� 		�p��{��]�%Y��5���>szo_�~�gt�u�?��Yki�4��9�}��ٿ�ۿ��j��'��6,'.X��P�WK�j&����|UV�ԥw3抜����$xq�m�{�k�Z7�&�eSm��T��ׅpЋ\6#u�^��4'�c�F���d��UC�$�!0%;�k��ţF�h��A�e�B2\g��:�d��Z�cy���\+~��	.M7
�8n�r�p���s���s����!�U|-���K��D��Q>�8�˵	t���6@�hR�{�ؓU��0K2)r�巰��9�K�=�ѨH;���Do���(5H}�Ƈ����E�B#LZh�v*�!� ��{H/��L��x�꤯��?��Q�!l�d��Y���(|��;#�ai~
��م����z�^��4��V��A��E�Ԅ+҅m��I���G0��A�\�ɗ@��<G�\ut�Z�F� �V���8z�Q��pyN���˿���������o{v ���҆�;��'�������=!͔��SG� _ C��L
79N�W�{`�#!�E%;x�֋�p�$fg&P,�Y�;EY?|�L���FD����1��C �x��'e* '�xKe�tKˋ
�qc�j@�RKel���A:�`
qS�E1e�
�~�x2F*�A�Ā�~�~�I//��9r�ڈtd�q�唔����Z�ܰ��&-(c �Q�J[�j�ښf�r������4V����-'E��h�Tj���.�ѡ��9�&0;3���o~��x��q,/��|�r��eT�dL,�os�Z b{yW8Y1���׸�X c��vs�fh�f��ZT�nn�&����	�?�jھe+֯_������~���_��/��٤�[�[Y\J����ɆC����
�9(��V?���_vQ#ŃF"Ӗ3O�/�|U��=y��rJ�J��������S>/r�2��$��N,s�(�P)2�ۥ�*�bw��NZn
ʙ� ���|.%��y�g��8�Uо��kSӦO�E�Oz��	�|���Ԝ����V�t��p��eM,�����ԣC��$��4>��&`��qp!u��mc��U��)�h֖��&8�"�(�������i��9�$����r��σLeC��l�*4|s�4@�G��s&������c�u&ګ�۠�B�)��\ɦ���� !;i���M�'1]ǐ�J�"�����D����`tN�o@C��hT5�F}
��R!�C�-�jUN��l�l��@7_f�9�3�\�H��oD ĥQ#��ד��/������������mv��䑿CZ$gB�~E�|~��$��t�g�ω]p�%��m���r����bu�182���ԯ=�^g�İ{<���p��}O@�&!����0՚r�}O�h��j�*�Ǹ��s���"î֏�LK���`9WE�B�)t�B>Ê�����JX-�9���MtsidӜ�39kSH���V	�@�j
��0~�(����@ȍ��O��Ki������#x�06>���)-��%�ó5I��/�D��D�wn��n���]����
�1����K�dԇ ��P�s*��r���K��S�����4vo�s��®Ꮏ����S���~8��h&�z�����{|u/�������̍?J�ZD8@��8�x��c#�1r�$V�f�}�t
>
�hx�I9o&���~$�0�u�}���Ζ�bp���T�KIf�̝���ԪĈl%p�)������f��Jу1|P�>*�
<.�))�E���@8�@_�7N��M�=Ѻ��4^G7ڋcc��A�Oc�r۷Ύ�x�R�8�T�!�� 2销�59��F�ɺ��O�}�Cx�soW5)���+�,�)��߾f�V�N{�����Ƃ#l4�e[�������LK{;���=j[�)/ǩ����y��wDu�j5�&۸U���ڣױ{�.�G�{����c��O��/��������Mzq%��G��T��0�վ}��=��|����������0���}~Vl.��bͯ��>J��}{�Bfi	�t
/��n��v�B�5ŢFc8v��|�9z<X�9}���@���"�w���_����xm�Q�6�GM��@���u����@F�@�#��*��+�Lh���%D͵���0����`�DSE�Oo�@6�ʩ��R�I�����9d��MK�\�#��9�,pM�(2�I�͑�~("ƈ`�\�kLbyM���a^�?�CD]	[����e�:��W|dٸ�������ظ@�o�k����CO@�BN�$���P��p���3o�K�|h�W��	�dS("^]YR��,]juj̴��3�8�`y��x��e �޹�L$�Z?6�%&�Ye��ӣ�6
v�ņm�4��m�[�ؖ��myN�8�Z[��J2�FC$1���L�¶%�. �6�l�2+�^=�W j�LL2���:j�J@��Iضž���׏BT;h�	�;;��C��Z��P	v� h&�C�b�.���i1ѓ��Q-JPK�L ��~��`����.�?�K'G,�ć��v�X7���,N�L��^��{~����Ǐb~1%�/�M�i,�*j1W�����a�ޛ�;�n�b}��g�]��ܙ�nj^Ꚁ,��q��M���q��ET�FQx�j!�,�^��7��{?u��!���|zS��x��c��Ǻ}�.ʕ��O_@�@�#�! 	�=rs�{�x�7�8y�fƱ4;�f1�H,,���A�vwch�z��=��	�=N
��R�_��Èv�c�杨4\�RH�{��?����/--`eyI�1)�B0�AV�fuZ.^��.�bj˨����
�oRvA?�z���XѼ�2�s�a�x�scMeҘ[XPU�DW��6�&ہBbi�����=��Ũp�Ǆ.k�bu!�)#��n��` W_}5>����jb��+]Ji'ϩ�g3��17-�*�?���v̠X��r����Ρe7/ˠp��@�)�M�nb�3��&	��;��F]��{����~�~^��u�D�?�O�o|�3��?Q��M��r*�����Q�ځiN�l��L�6��_
�s���.������>9[$�eN�<˪xn��r.�B:�{�K�fn~��8zz��+qqr
3��!�Uh��C�K�T�oN2Q������������UC1�P�ʏ�hT��Xy $�ݚ*��7[�A^��Gr7���M���]�]2,����-�v0k�߶�t��.�c\�8��`$�&�@EN� ;b4,�KpSxo5L"�P铏J��JC&pԄPy����n>kD�|l����D̊���]-��(��'�y��A���^NWH�`�t;�$0&�b�̸?��&��h��h�5�׃��073��Q�Zt��P���6���7S���Q>n���~��� ���)�7ު�CFe��"�8ä$���Q�U���'�~�jS8��|L~/?���IĶ{Y>�a��v��]sD��Y�P5��h. m[��G�3����f�'c��LPc�|�Q1�|���51�E�P�n�
��k��Ҵ�XH�n�
��w]���G@�����
u�卡H�j��p?�=�Ĭ]��>�K��RN ���7]:SB�"^��gq��Q�N�;�ƛ^�*�����ȃ?�ٓ�T�o��\�F�s�.�b�☦���E�=s�([X^-"�1�[���=�a)]D��A��ڒ���3@���΍:�|�:z{�8r�1\����7 m%�} ����?�я���TȨ��|�S�L����5Q���)�p��Ed�uT�ӱϟ��[��-d�f0=9��G�Q�j�&򣯻��eM��5�H��cGpij� �ifC{�0
�,�7m݁���h4D�A�P0_AjzGqNǃ��,-.H�k�)F�bV�����0���8δk@�b�f��U!M<�x��c��f􍛑eTx�R�a���|�I��j�PԤ��@o�Q�����:@��N�0A��5P�����F��UO����=�9zm��Č-��bZ��S9m2�4(�㈸zm�=����T�h��9�٬lem�ϟ������N�Y �m��:�&2��,�-��w�1>*7�t�~��@�]{��s?�'��g>�7JӦ��
�C*�״�F�5N�r� ��aVƣs������;�w�^}��W��E�h�����#�V��	_�+Q�6%�Y����4���P��دI�T��X�Û6aznQ�J��	^53a���]ɸ�J8D[�&r�4��.�͖��r-�m�
��V�����T���TȰ���_!4��QH��I�f��    IDAT�ľS���2!?�
�"��쬭��y~���������_�g��2P����53Ȋ��Ku0��%��p�{��B�.+R���?�@X	���y��w�[$pT���f����]`����O}Z��̹�X^Y�������պy�F�����F�M]��\��' ��������G���s�)�tcnf�0�v���0PMH6Ԟ"8ݾc^����G�ɓ'�{���n�M�e���ZL�e�������xd�Z�a�{l�(���#�R�m�2[?����K�b5,�y�L+��m/ ��c��=��B�j��n�y�v=R�C�@�����H(� 8Y%�dt�~��׌�A�fSg���µ�B.�;����
Y�(��^ �W�7�7�>�	L��z)ح� T�s�c�F��T�H�#?��ip��̟
�N/�&^p�-����O>� �������Y���e�pCx��_��cjQ�(����^5�2.f�W121�ZՇH�0����#[����*��D�k�[x��Q�����@oB����1Ը��� *�{���=@��Bzs��x�S��r�V0�JH�x��%�st��k,�\�#BWZW��*.�>�s�A��,mG�����̫v�ځx(�
�I6_���$B��n�t	�B�x��	oV�7v`h�vT�^k4���#͡�ύ�r2V�Шs���޳Z�&+�Oҽ��&���J��i��4��<Hnx��h�Z�Q��
�t$.oBm����H����^�F,LVLJ�bZ?|�`�S?��*�t��Z�J�|;��\��ً���������nG�4�O�N�:�B�����\��������lOۚ>��o)aT,���:�ϛ�z/����Ӷo��|�ae�e#�6BCj
�mۢ�����ԛ޺i#�]�_�������/���9>JZ]aeŒ�+	�TI9B�a�%����lƜ�a����r���%DV�!�;ʣ��(F� � �M#@R����Cشi#��;U�p�����&0���\����U�8�J��ۣ�B<䗠�:%���G�aa��eLL�JlI_ ��/VҤ��S�s%�u~N��� zz�.;�*
�p���f�l�ۙ������^۾�r�Y�c��f��ǳ�r����ͤ����J�6�bd�n��,4b�c>�f�4��Y!��4!��}���4z��������3��l&�����~��߆�� ;@Ŀ���{��~i~x�O�=+�z���ʾGS�=s^��nc�u�}������k��U��}�[_���4��R�)ܖ�ף��V';l,�8���&yի^��|�#x��?�o}�[zx��رG�>�q�C&-P�`���ⸯ�����}����0G�v��[E[H<��U��A�ԏ���~�\8��-|��>���W���V�&Όy��[M�t?
b�4.��ޫ u,)��u�{(�ok���$�kFg��b^�e��cϵȖ!��
�Qi�PC���\���,ƃ�H���@YZ� ::�����ZY{p}�
��2�.`��	��Bgzj��߃MÃ�1:rNk���֨u(��?�|�$�
��O&�q�V<}�?�RՅ\��kn�[v^��U�Sd��{� ���|�Qak�Ṱ�#������4���A� j�;>�G~׳�Q�Lo�z�<zf�m-܏P����Μ�@*��|�24Ѭ����]���\8s��1c>4kED̵�`��uؼq�;���X^͈�nz������+�f����Jj	��n�mB�E�F�Bg[��9�)�^^��ʂjҖ�9Q�c¤Za�9)t�xXіP�,��
5*dX�ܼx͚G"�iP��t�opnƋ����F6��d3Jw�� zZ��)1��9܆T�Z��i�1mDl�����t�I���:d9Nv�bP�n�Ȥ�)N#���.��˲�7�6g<�i�mJ{H���)���kq6cgӐ@�m��vS���y�	 ��l(l���Inx<�xï߰N�g����6��ǟ�OH�9�5�
4�"TKP���aU,# �WT2�ż���Q'��:"��*u�q�R��)R�-4���j!����/���vnǫ�{�F���:{:�'��������̜���&���*�*P�T�:�(:�QD#A���LOH�PaK����������x�|G8v;>:���i,���Q)+�Ɠ�J�gEʃ��,�J�J��i;����v c+\K�{ȭ=��Q��e��w*q2Qf]��X�i��k��F"aZ�Sc2==�o�;���C$C�V�M�Ʈ������.�������w�L�K$G]���MJ ��ۏt����o~����=�yV�YlٲUbk�3R�|��ڋZs�`Xk�q�f�Y-"�;�m��_�
����~K3ڏ�>M/(>g�sӳ3Zs�P����X8���l�K^������S��æM����C����V͚#dv�ZȨ����X�dX;	�w�gvoh����S,���J֮��BFm��ߣ��c���RI�55h4Z�Ə��ѣG�s�Z����)(mxݵ�y������h��"A-�am��%�b5*�j������T����!��}h�;Qi�-�UX�}-�-97��0q8_���#�t�կ�v��bJ:|M~�?�:}�N?��nl�ƞm[�¼��YI��$,߼e;b�N�$��0�dm����|2�|���Ï=���o Shbtb�����{^��T%z����#,PQ�L�.���3��܃F�Q!��U!w}~�P����C�|v �~���[�>;���@��M5�=?��J�;��VU�lv��<sK3��4
J���<�|�CwW��ne�ԛȬ�Mn̯�S0��[v!�P���<|�����wxeWs�:�fJX�5��DPg~�|NrqM/ͩ"�[�9�J�mZ�YtC��c4**����J�Bsn윇����ˆ��z��
ь� VZ��9���H$,�����fgTI��c�Iy�֋�Ia6�X7�&�P鈆ѝ�	��NO�u�PO�Ԇ�����r�������k;v��AEq�G$���U�OcX�"o�RI���c��h�d����ѻ�VQb)��͊(� pc2_XE����������M���~nVŤ�0*�#,�l�YA�&l��O�C��
d�j����e��i�r�]��頨��5x��E3 ������z^t�=��������Zh˩4�� �oބ��9=g�WWWE9�}n��}/����_�W�D<���"R+��슋u sBF����:Ӳ�S-�ܙ�x��'p��cXYM#�-�ˈ!���ׁ"��d��2���[{�-X���nɶx��C�C�2,��]C��]j���e;�*�P]�pn��af��W��S��w�G�<-��^���J�3�oX����t��NM��Z���Rk)j�X0��Q�C0���^�h��_��� u?~�'�=Z��r4��C�yۦ���8q |�vnߊ���r+��Cb��9y6u%(W���64 ��}�,�_yͫq�M7;�c8v��a<��S���Ta�ʛ�?�LKЀ�mS|�[o��{�-B������6����[��Ѧec�הm��';D7Z���^���������_ ��em�/���0Դc/3*�0�1-�@���}�fg�ٸ���s�~���<q�~��$�?���an�@i��)�fL{.G����ތt��t�	Ĕ���@"�F��ő�~�|vqa7vm]��o��LcG��4�ťY�ooظ[��@oϐ�����B)�#�U���;1>1�?���`~%����������Rӏ�t5G�����Q�h�-P��w���`d�"8�ȩioP�۵���������g����Jq]�zӱ�3�y#AW�aTr��F&SA�L��'�O�������ɧPZ�A$��.�aN�Tq�K�Eoo�n�H<���%�3yLLN���� jM/:��Ȯ���p7�aC��m�A�8^��~� �����-6��R8��4���9iL,Hq���f�%��{���J�b�i[P���,@_�d��	D¦�M��C�@�Y3�@P7\<W�=�PS�j�5y�9oߒ���MjTl��ҙ]k@�X��ۙ�������*|�,"5^�*����>^'�����fUjiٽ{�頢3-�7?o��YEX��<�@�02^���=����Ӛ����@�~�ҧ���3Xf�TW�E��I�3�}��6`k�|�f���5��qf*潬$B��Mf��,W(8fUm�U�)�-���;�/�(kU��Q'��ȼ���.�{T73YzyU[F|Ib����Zw���pݵ���	���Z������opX'���xͦ.��eă~�t�5ȧW05>"����� fqx�:�yy2p#��~������+j�8x� �����X!k0��b�[���0�a��:���BLk{�m����q���dD���)��T��u�!/�႙�f�zð��(ꯆ6m����x�;4�ª;�+�X��ĀG��7���ӄ0[��6m6-��Y�ɠh��낀����~�zPk͍�[�	(=��#z��n�!�byF� f;�-}\-g��3s(�`��h���z�����Ǐp��3��m\?�{�bRޛ����Ϳ�ƛ�ַ�w����X������bI�����NNL;i��� P1�Z5�\,��K��m�eJ-@������%u���Ҕ�#Tms�����5��LV�@��Ո�#*��/_��%��;��9��[��v�#�����g�GbZ2��y�S���0{l`n�Q�W�*�� ��T�IT���
#�m"5s#'�:	.���ի-���㚛�@0чg�9z^bޏ��;����'~�=x\y�t�1��m7���k��ȹ�`K�Q���I�c]����<z�zE �x����s�s��m��}����#���� Wv�/-��nL.��ru�D|��#̳�ӱ����7��K����piD�
b�Q�۽�����w�����;ӎL���|��c��ƺ��Pwy��*�i,-SX���ӤheG�|+�h�S����jؾm3�x���}��I�NS9�8�:�i�Vm�t	�l]��:"�㎛��D�`?F���1>WA�B:W��#�����s�<Kw�%�%Ɛ��@$���u*[B�1 bU���fUm���,��HX'�@��*\��J��.mh��O�n���(�M\,Q(��7d�"Mň��T� �Օ��F��%EX>wa��l
=ɸ^}j��Ln��WA�&�i�,
�^��x�[J�(����Ҋi�
J�����Y�)��'���%��<TH%��k[}����6?2�Ċi-�igf�fH�Cm�<*�q�q �˰^�Ǆ�0������<���$�,�i
4�.�[�X���?���CAab��MȜ�� �׉��]���ˠ׏��>�jl�=w>O9�s��j�Q?CMӜ=�fWP,��4G�iuݨ"���;���ɉT+t$�I�\������ܙSX]^|�o�6����,&��ojwx�>�����_����/TL���R���Ѻ�����mߴ���j��_��R��t �tS�Z&��N�-�-\�6L�e��+��:��~��ذ���A���������r��k�,�R��VKu���q\�O��^�d��豤�[��Ԫp"��}-�^ģf�'b1�K���;==��?�tz(��j���#���jp�uk��љ��}��P�Џ���8s�8�A::b�ʐ����sg��ʖ}��Kyɽ/���[	��|����T*�1�ӧΫUB%�b�ε�$Ӻeت��L���W^���!0���y�����O{�:O_	hm���>��4\ܷo6m٬��$���CM�--��Ŏ7+#��
����B���2�5�tc���B�N��c<����=������hoT����n��1*Uw��0�$ʈ�>?����ɷQ�<JnQ-������}��zl�{=���`Nm[2g��z1}�(�|�@Q7vn���d��>R�]�_�
�B���n����h�wtu:���Hw_���p����>��TUq��Æ�pn|���pI�i(�4je�vձq� �x�A\�F��B�qy�s{��?����3w�\n��ٿ�f�o������_.U+��|���x�=AW0��ۇ�L��Oai%��
�}D�sSp���V��(��T�q�_��S�`����z�᧰4_���Z�&�o� 3�#O=��J7�ۇ훆p�Wa`��D� �o ��i
=q�j@�'�PSt�p��a��������%������E4�-�:���ԩȴʤ��_��G7Y�zI&u���T��=�ղX�PT�E�м19Ya,�M�M��V�7y�ZS�*������� -�a�\���(dVŨDP�czzjm$Xs� ��jL�l�I��ζ 7(VUf�(�giqY�K��ǭ�O���$v��휕�egJǀ{���l;�k[Q��lR���-P1�]' �i�EH��Zrޗ��U|?9���N�14.Y����%TE�T���1�"�&J^㈎ˮ�$i�Ն�'=/t+�R�U����)M�BӖU�hO�e/~:�1�BA�t$%¦�fie]=����ɳ���xc�3r�����Q��;�����+9|�o?W����^�+�Ҹa�~�>sR��l������FS�rWo�p��S��8:���e��%�%d(�u���Z����6�~]y��Zv}���+q|�+��C�N�p��i�~MQE�!���ٳ��?������w��?��?�ŋcغc'J��fLMi�u��vZ��+)B��۱��yr��͙g�& |(���`��#�h�yg�Utݙ��{�q4�S��g�Z^�A|&��ػK�!����hwoߊ��p��	�>u\���}]�+���b9��s����59_d^�W�/�Wm1MѺ�B�����XYY]*de�d�戥ہ�֌|x�$�/bL�<1��zV��&�u�v0j��L	����@Ȋi	TȨPg�a��5�����|�;*t���"ѯڸ]��?�	�Q!{]-�T��" ���S�o�������D�q	�[����\N�l��n�G� Ax"dT�Pu�5BmJ e�9�(�#'��͞V�׀�A�;�p�w"���^@�?��7�ĩ#8v�A���H��+�\z�]=b��z$�g���̔��N�:�f�#.e�����<G�?��z��݋��Y?}Afo����~��3+YX7�芅����Y�>��,,�<���������j�Q1��AW����>�g	P_*�7>>�w�;��TV�5����M$�aD|-�z�I�;��SD]��""����}�(��d
���.c+E̯,�����9�����Al��]w݆Mۆ���1��=�������.W�ly%`�9[2�P=w
��cb�?� ��:��Nt�� Oaf�m��O�-O÷Z�0*M��>�
��a6u!w&�G&�7"���Q�;���wx��ژ1đ:k�$�A��n��� �r�eM��tĕ151�P�XgS(��R���v����NP�՟<��������KNl{�T�Ĵ���`'wVWWL�ò�Mg��_����ˉ%q<Ԯq��.�Δ�����n��%����AUΙ1fK���&�N�猭�$$I�M4E�dF,P�aѕ@�`Ql�eX$�5�:�(.�y�{���&3��n��J�����_S?�BɄ�ii�Ǳ{ꊘ����"��#��kC�d���;�~��7�Q��/��ЬU�?Љ��*�n��:��EU�oy����7��F�y����g��cO�칋b�%�6*H���}�ב�������{]-�n���ڵ��ZGk���Ƿz��C�?����Q�qBΏH0�x"�l6�1u���[����&>��O�gN��k���ONKL�{�^k�ʤϒR�W�j��d;�����\K4�_1s.h�R���ݣuH!����9�uV�k)�ds�	�Īx��Vc��Ȩ2��� �Bt$"�gV��0�d�Q�~    IDAT�ZO��X����>��LQ�+_�J����*�Q"�#�$�B�i2*��^�F��ψQq���l�aX{�-Xm��_ɰ��6�Kc��o��G* .�^̂3�=�w�,�^i=�t�-ؿ�
-\4#��W�����z�b;��Mf�l8��� �MT�*t�����x���Dnx�:��@(��TS��j�E9]Ð�BQ-���n�j��l% ���KL�VS�S�Y,O���3������=Ս�=Q���p�����c5��s��J�3��؉C8�IDU��6��0PȦ�i�zM�qH��<�ZE�v�^}8��K�f]y ��QN��]�ds�8>���ev*���N�ۺW[&?`RWڕ�����f�5z��04�-�ri�>*N��/�=C��ȇ~����\Z���799�Aw�3��E������Y,�P.��6�*\8u��4��4���z1LC�M�رs�6�)&�CRA�i��@���� Ώ�W���j~��B�J�p����׉���1��`|1�R+��.�+
?Mۚ�r+8~�	̏� ��*�88���#�9�ξur�u1\�1Ņ5�~2��z�~jE��u��1������ӥ��Z��M����س�~jF<2S���on�{����ˤK�mV�ר� (�#��������n�'��L#ٕԆ�C��N:��d�d�W�7��M����}]���~m+�i����i���[��oT���5��1ɚ�iP�� ,�˟S�3�~XY\dZU�����erHx3���H H��*�yG��cT�)��y���Ej�P��Jg�q�lk�Dz�|΄����V�ҳH �1d�z=�YӞ����׀?�S��BY��*�+m1�L6%�C"ىL�$�2�aW���]�GO�JI���=�{Z��Sۇ�*��]�O>���-[6�mo;���7�����N���8t���dځ�L����h��@j%fB���Z��-�������3��~���~�]	T�ꡰā�BN�.���'�s�^<�Џ��\l����g�_���r�4©>
�5�fZ�!i?�MS��4ܽ{��Ž��������P��%�EZ_�&L���%���Qא�53	dܪ9dZ��P�S��i"�^F4�S�G����P�z���$�
G4�C�E�+_�rY+��>���C=���E�ы:�FFF���`��۴s/�\��m��W^ӟ����*�)5�ާ6�c�2��'���/������[q�u���4xd*�׾�5��y$��Ԝ�A35I&Mڶ�aVk��ᐜwݝj�)`�N<G����W �S4����������J��;4_lv�Q�j�5�h�3;}�N����7�7=[w�C�PB�°S��0��ة�8}�Q����ҏ{n��y�VMQx�M7+1z~qA�w<�9J�>}��
�����4\'�F[&�|O�>�\���L$p�s��d��ruT���j!�/]��y )����|T�x�'bTT��u����������� *c��\9�棧/��/ޓ�aL��G�PǥKHe�X^Jk*�YN��?���Y��)��ԋ�}^�����]�]�[Z����?�����_��(��'�8�cϜ��A�jo˃��A��Q�M$5�=�ZƩ�l؋�-Wa1E�k@-W�����p��㨦�
�F�m�C�u"�;�-怰��T,�b[?�QqQ�Fz�Ŕ֠�K���ހ���4�nf�-UD�̪�w��F�;@E0�@�ؒ�9ŕ*dTTB^8@e��e!li_�7P��Q)9/qU!��%�4�F��#�h$��N
)���B ��AWP��@��kD�Mm|vԑ��y?C�8mK��r\l��m�}�Ǔ�����YC[��Z+�T~f��� �0�kfv� ��A��[�B�s�l�k��	c�&�"�� ��!�q�E�dh�E��1⍬�c���ҏ�t�R�]�f�y�0^��{p���8s�<�o��͛Q�5q��1?y3�b�JyN�q�\l� u���W}����N(����?uP��,��x����׾�q��H�?�c�N`rj�3�ȗ9�k�	h�nY��kwe%m_��+u
�1����q"���[Փ�TX�&�Q�dT���E�DȁO�]y��'�78$q<ǆ	T���0��d_->x�s7��	��x4*��Ƕ ��F�<�,�-0mF�5b[�V٦�:��7
�N��(�z�>$����NK��)#��+�r���=
U�x��!�� P��i�׼�5x��^�Te6+�{���lvzV�S�K�#�"�V�z̽�k�cڎ����� ò.���v�ݸ������c9��,j;8�=�=D�jTG��n��&�T���R�w��]|�+�(Q1�k��]2�k�(�fñ9h�F�"L_ϕ��f�Ԫ�'��ܰE��D��:08�}si5�ӧO�Z)���K-�k���b�2o�~�'7|*ܽy��\5pcz��gm���a�z�]'�1��$a,#[j�2z⨥�q�'߁��Fo܃���anrGBOw��#6l�$V�R-���W�Y>�G��C҂��IMu&;{q��������_�R&�L��`g?n}���tI�R��Y� ��'��Yӄ��f�f}�q:������� ?�s{�u|�?���>+4**��돝��{�Xo���?�����r��l�hb�Qg`a�$P\Py�k_���{����U�r:����7�'L2p0�G~uUoA'N�@�R�fU��$t��V�w!U�a|.�3�f�i�>oك�|M!d�L=�2�ϟ�i���D_qdS����:�5�Ѯ~�[��T��Rέ�iT(�u5�j���6�MY�3f�&7��/hYg�fe�E�S11">_�����ޥF���L���:}!L�@Ŧ'3��R*�O����TI����v)��e/{n��9���/7,����%LLL��mu%����_ T���X1}a	z��B��e78:�����`���$1�����d�>4>�j����^�-[����K��o|���~$�cuOu�xel���~�O�,��ڢf�aPd��ބ�D��Rdů��Jm&�l�T͖B��F!��~>^��;���Ilݼ���_ǉgN��`���_�Ξ1�1��K��S���jV�q1��%�
�
'�b��9E��`�����}��w��>�3�/Mȡ��gΈ��_XF����2R����͵��o'd�Uտh-��~�Ǖ@E!'	�&b,�i���af|t���ҁ��I�j,�c���;��G?�Q�'���C���E} (��?�ݔ/3Mf�ô�Pw��97ΑN
v�G���RH���3�v|�&�L��z����u;.�.���Ðbo�%0�}�����׍��<�>��ފ��Y�NO�w�8��q_��'m��u��>$s�i}<��Ø����@� gl�|��
[)*P�7�E�hG�A�eT�>Y1�(����q�����vm�/ˀ#5qؔΏ��@�EVwW��
��|_���cddD�"���5NnL�ȨH�҄)pP��@S+�^!襠u�����_B�����xg�D��F�O��=-�����Kɨ�B��F�KNr��$��X��F9/�)]��h��7lA��F,��ĉŊ�.A�p��!3�@�y�]x��7��S���)��?��ە�Mc<����H�K2�㹚˗Q��1����\��jHl���߅Z+�t��b�8v�u�����^2�L�|����8�|\@�*�Ac��k��v�K~�O��;��i��ʕ��/����bZ�b#r��S��F{*u��l�/Lcn1�/,��S�c��1L�A+���Q��u��k^y��hY}�n�K_�w�9?����%b�8��T�\��ܼ4�ᆇ���bfv�V ��
3u��E��f�۶�0+��@$ d�'p��a�M�G��X���@��&��	��&咦\V�B�BF�Z�3�`�E���hU9��BPUSL�[.VuI���J�;g��7Z(��v
+Օ�d��ĵdTT4xh˹��рGf�t%�Ȧ�z�4<#=ɞ4��뵢Du������-�u�=JO�Z.�0?��.�?��|�If̘�Q�M��޳=HLuRS{��o5V�o5v4�V��W�|�bJ!o`j$��,;7Aܠl �4�r��}��k�ݧ��3�����'����_�;�A����a���RK��T�E!Pa�Ea�K���2�S�M�SBƃ��U�N+�#�xɨ��JZᗬl�9��;���=��g�/��.�a?����H������7���ҳ�j�b^�mn:-���^�~�ʤm_��L��i̟�r��g����0�}�K9֦��ع�p�N�<��KX\ZE�B�7C'������v��J����v������0e?�2���9��RV�B��>um�����2�����="'֧O<�5L�� ��kG�	�F��x3C�7�w܄7Z���T���{��D]Ų@6��ցt�(q�T�wZ�os��a�l)G��b(@�`X��Q Cs�PbPE�GeK���]��Gju	���]/�[�fN��������:��e�CQo˅Gy�F/i�ultR���51-�@E�èXG�v�i׈Ƹ��&�-^{O�A���zIc��I<�\�_�:�|��"�i�-�,������=����/��ٳb����%�
)�~a�������/]�m��Q	��41.�}���n��V1,�+��~%W]{��J��G�ۍ�')�B/��D�ԫ���(T��Æ�����6dO1G��Fٛ&b{���>��G�Ne�p��;����)|���C����}�w%�7Џ�ǟ�k۵u�Z�3�H&:p~d�b>��<2�

�
��2�	F1�i;v^}=V�U4�a4>�������4M��7�7i�A�r��eF���T�b�����o�5@�P=p���xc�F5b��o���qLϭ*�G�7�2fF���㏡�:���ox�+��7ݏ������~���G������[U��!0!U��^э�j�Ϳ��q��q��N#Wvctb��Ex��u���h�:��ŬLk\�,�Ο���IT��#)�Q��7"�9�'���嗠�2i�+҇�����5��c��[j�X4,�]*�Gŀn,
�4�������2���R����e�
����22l����Eq�#F%�^����T"EFeiI�.4�(�)�<�%��.C�sk4DR��o~<%��.͓�hD����*ܴxÚ*���!�ѐ��'`��蟡�}tQ-k<���PX"���M��ֈ���x#��bޛlܴ���FT����j\��W��������W��\ވ�������vL�YMfP��)K��QdN>Q3dĸ����I�BzW����S*v&X��"8��@/��_�{_p�'q��{��~���u7݌��y7������sH�3
��H,��k����}|<��ѡ��B!��EfwTu�v�خ��W���<z�(W����9}�.!�+�S��:����\-���>*L���1�p�_��@E@�mM��R|	9��D�1`c�i�ָ��(�ż2z���w���O�'��x2��y��K$�"+��קI�LN�,c�M�[�3w�>�`Q���7 @GXO��gU���=����Ű=�`;�����ȫu<�M��T��yN��oǱB�pY`�.����2� �� �V�e��}�zM^���:����sd '�rx�~%fs�a ��ёQ��''f���]���d�s���A�AmYL�c�6����ǭ��.q��5�ǿy�+�*v�����L���"]�ј�o��V�x��|<�Ql�}�_��3�L.��"Y
�M!�]�oFa�è(p1�x�C�w�^�f��p4*��t:��C�E5��⧏�1"�=���s��Quu���*ިX���R��ǋrZ����Dv���|.c�4 ��UA"�rsx��!�<�d����ٍMCØ���s�{�����qĒ	,./�%������%9�s�t5U��j�J-w �Z�P*�ڈ-�����m�\� M��
4EB�p_���\��@o�U��UCOO�|F/�����bTv%>����s�
�rq>�[nFx��3��'h�V�4��41>���4j���|�����(fF�`i��"��M}x�K_w����%�$fsEB1t������e*���9�[?�Tj���ضs^��{����q��SX-4Q��0�T|Q�r�=
X�'�͂o,���gǱ<7FlS��?�>g�6/"���Kɟ�êՇ� J�>*Ŕ*uNQ/A4S��k�G�b=�����H-[V�==��x�PP����I����JH(A�����j�T.]*��IW�)���wK���h�
�3]e��ъ�v�mx�[�"f�π�*+T��$���׿��7W� x�ѐ{(8a�*U@�߂X"e�;9��,?�
�4���b�l���y�:����1?���N�����l$����ݽG��[�����	��_�9����T.+?��JY����U�[:<D�}a�U�TSd������ 2=�8�IP�נ׹v�U��qD�BZ^�J6���$~��aǖ�:hI]�9{��{/:��p���NL"�ex"sg��
��NB��.9�ɐH�ZQ����pB��ͪ��W�-��fM5�-.�ob~~Q mfv^�4����ȡؔ��R��p��ՙ�k��_�]�8��� r��=����U!��A��qj��&È|~�XTN��vluvv������xi�RG(5���~|(���Ҕ�6,5`�>S5����F��aҙH�� �:��(�)`�S�TT ��Z����B�Ta�9����gr�C�9�z|A�����$y�ԴeEP��Ĝ�0ɧ�n��|����q"����ߺ}�l���~Y��Rop\��k?2r����&3�v	���t2����iӖآ�{��i��n��������x��]�-g�JŐ�D��/�w�$��yǶ��f�>tuw(ٙ���}s�ٺ��d&�ۃ�'���� ѿ=n�N�0'n��t�唔�hB�P"6�j��z����4�s��q�o��v��!��ܚ4-�p�{Qs�Q%�d��&�M7�� 4��<W�#�H�up�9���_A�n���b������c?s�F_�Z	~��]Yg5J$;;��o܀�u�0;5���4jM�c��9�O�![��Pㄗ�H�w]�;���#S���	�ؒ;n�SVz25**Ү�˚ ��㑇��ӓ(s�3j�������>�z������J+���G�~4ҽ.�@tO��4:���,���̙���.�aq�$f�O���G<��t&t��jO$:�i�Vkr%��U#���FE�����܅�L-�P�����cv1��;q��[Pmy�-R;BD[�x'E@��Yd��Ć�Zm���
�#6���/=sA�Mj�
S�˅���a�2�f�k���V��I΍�M�Q���֡��G���\AcqD����z��2�H��$�m2�ޤ{<-�����˝�+�@O�63���>2����������_�J�;�5]*�醉�iL�O�F?t�)�j5����mK�����'mB΁�������rdL���9*NEf�2�5�C�B�E0z58F��y/� V;��1c����^s�a��ݢ�n�l4�������݃�~�s��O��Պ�F� ��^��SZ��M��!k=p`|Z2���E��Z�s:�H�
}>�'j�D�P�f�dl�׍Rj]]�G&��Ƶ�~�f��A��˫� ��e�Z�{.�u�Aʫ�p(�D2*�::zA@/bF�KUwg6��J:�<�L.�d�Ӭon�p�ɒ�<�,(�u�FL���T:��2.k'���γklo�����=��Q��SM��4����ڮ7�n4f������F�K���B�\tB�!��^�ؕ�~����
�k�&j�I0���K�����=�2�=��.���x�rkH��b|Nyqa��1q����TM    IDATz|uS���L�_%@��ټG4x�1���S�hVr2��f�Q�=�=�@�	T^���{�A�wkLOL�!s���$Ƶ��W�/�!	=�@Eסe։m�XfTzN!w%Pm_�~i%�A�g�F�>�q�m$��δ`;�р�L(-M��� x!��靦q�Ծ��Of��P-Ž�N�M.fK��F�6oڪÝ��������}�����`��]*d�'�015)p��:������K�Bh{����!_-�� q,:�7��ׅ,����y�s$�Y�%�P�
"�B�ʙe��:����t��#�Fh����3F��RW/��s��XE�T�6^�F�ϏM*V�L ѷ��E��z��nMya��xF��t�O�R9'amo�).M���r)*D�����]�����3�
FE@�yݑ���O�w��<]�V0r~
KyxIi6x�U��-����㘹x�jN�LJ�C��iw���/�6G8I������(uv F��cS�[�������:����!�ѫ7�Xk�EҬѣPm�w�,��rӢp�����M�/,q��h�ր����T8�L�B�@7�[?��\|h!��a���6R���M���~��KcX�_��];��@A�㬰�}�0�X�:7iS������A�>g)�*�¬�s�3�20�����D!P��?�k�]'kiC��S�Q��w���G�J<�M���gn�V�.�æ��W��M�$:[7��:��J�}ͶM�<=jh������q��Y��WS�3"<3�ȱkZ|?���"뇆��t*Y#>�?�|�+���\�/B��kǖ A�i��J[�QA�>0m������׬�Ή
��g-���K��;��
W��L%�:7��>� ʃ1 ���ja���XXZ1����P��b�
GO�*]q�(#ςS+�m�@ᶫ��:��J����
7�$����Fo�p��q�@ک�vvdM�T�WjR����vPPQ���40��
��u��h�v���	���;�	�X��TkfR'�8�xTx�	0�sX�5dW�z&S
t�W+�%�Q��P.�V���B�j��@�è�BgJ� �2Z'��ޠ��0�GŁ�GKSkf���b�)�.eV�nUy�I��Y���L�6�Y	�x<��\��N�f�z�d���oټC���T��!FLkD�<��>&�#�V(��곀�2����"���7�7r���6��� 1@ο�ζI���!8ZY�hp]L��R���$��Q���5����ic���4�I�7��X/z��t�՗�]��"�^<���؉��a\����Ei�����y�f�p����Y�"S��;܏bÃ2Y8��5
{��"Z�͆1�@���@�'��ԧ��QN�+�E�����y�;q��B��[�p 	V�Ѱ������X$j��!D���0:���΁.��D��ݏ���h�#H�J��-����v�B���zt<�r�����`�Z?#�FPn����0A-7w���O�����h�����N����V0!����������I,,e�t�R��G�[E����Ӈ1z�8���;T�@'Fc��qy�0�1����"X�xt��ڸy�{��p~t����"]hbz1_�][�����GQ�C#ˢ��WS�]���<�+����ц�6���ʪѼzL���]�"�<+�}�'��N�bEMZ���
<��mڨhlt|-{&��KC��6_(b��]
��hk�a��:��sL}�s�a��JL�11ƀ{�'CT)#�q��cc(���`n�.�� ��}���w� ���L�����q����[%Un6�Z?-���A�I+��i��j�V����I(���ی=�,�v;^l��6G�h&OH�M�v	����P��100��mԷ�~�Fڿ�_�W�Ͽ�"�.��P/S(�O�ZVr��H�����Q!��}��/������L�wBV��9��$�U�j�Z%��rl����|%�5M�67S���cêmh�9�rc�t;=.>��j�4ɨ0�#T����ł $�'?[��!r�=�soe�y�y>w�o�T�eY��$gwB'N��q�@�i��p��L�24�4�!��n��%H��$��x�,ɒ%۲�����������+U<̡Ϝ�9.YRխ[��~��<��p���3	:�%ז�'NL���H���v����~���;k]��[������uE���+녵ӄpX#��)�)N��q��!�S8��9�@�(��Q�V��������&�=��q|��y�o��*���{��du�$�"�� �|?lo�O�����9i��e8�#���*]Y�)2�$xo-�4��G�V-Y�^'����E����+{�{�dҸDwU�����{bm\w�M*����Z�Ba<{�8��/�|���iힾL������%|�9��`��rN�?�����*�\�
���QR�3MC�n	��������֚
y��?.��V�e�|A�}��:��p�Wn`@F���Kjbs���WW�[�"���m�F�.�Tm���Nr�"�1���֦�b�c�z�Th ���e3I��R�0;c�z]�#���(�KǺ6��Yui�^8��-�=n�XG�'�j4њ M��q7�[,���QL|�d�C�68�ٶ_u���CV��l	D	�8��D���"�]q5�18c�;�+�q�*��ջ=����(T��2����Ͻ2ȴ*�H���ǧ~��Oc��ʦlf�m/��=��%����kW,��Z"Ұ��ى�men�:ͪ
��4���%��֭۶�-�MHv'��vW������s��-���jG���;����M�g���Z$��^��ͼ�k��¬--�Y��ԁԣP���:Y�^��{]KF�j!}�f��)+/�(=��e2׳n�H�8��L������R��N�� �jw��e��y�����)9HEPd�l��H&���mcC�u��S��l�Oɖ��L�i����]ួW�C=dozӛ�i�*{����ivnA]#!�A`uL�
����R[���]�ҭ_���K ���_�� ��pC���<���Rl �n)(zB�ؤ��y��q�g��!������=m�z�)�$]�����RiaAY.!�{�����Bg��du�N�&��N�^����2�Q�cK�sv��KB �)�*����61>nW��m�sv��%���N�#B�0������mܤk_'w���ӕB�D�q_.��B����I���E(���Թ5�a5-?PHޞ>�5�q^����>]�����c����k��P�"-~�;�*�)��ё����Q������P�\	��USFq�՛5O��ߡ��Y��K�Bť��a�Aqρ��$5.۱c��g�ʊ�*
E�k��UR�������q�I�O���gϪh���B$}���N�_2�\'м<�@�L���n�Ŀj�+U'c=ۻ{�U+%���h��H����J���Xst��s$ʟO�@C��s��B����@�0�e�ћ#��N��~�6,L�����Fb�^��=yo�1a���ە�g}��ȕ六Q�&^�8��0���E��U h?�Q&�/�E%��R��=���6c? [<��!xT|������x�}
#�^�[�7��*����.�j#�BŒ�ִ���yc��/v+TX=���mx0/��t���%�g7	$�4�۴\�o�H˖�/؅�Glaꂔ�jI�H�
7��\����){�]��]��m��.��a�#��MY4��zr-���9���9�#rvǩ9��S
�M�G���'���cV�L�H�*����o��Ͼr
K�?���oU{��PI��R�N����K��3�>H�|ҬR��S/>ggN�^�j�ʪ`��6��x����f�1 ���Ge�uijΒ����,����y��������j+e8qk����ڄ��z������8/TE�9�uy��Id�pͳrЎ'�@�I�W.[iq�:��E��cz*��� �B�K%c�}�V���8�+j��/�ɭ�
ț:x�Y+W�:�!���H���:�|��[�46b�]�G#,�;,�S'N�5�NB*�^
�V�	\l���CC655#�����U�D�l߳0*�1�_R��J�cq����l��q�+�<�l�2�zb�6B���s�t��8���t"o4T� ���NX�J"l"e�FG�C:������k������+}�i������6�e�n����S6;}ɞ������6X�|k\O�@�vۖ��llx���ZR�����������d�!g
(������ӦDэ!*2]����Ϻ�~�o�=���:r$��9�aB��kȳ�5f�����e�釣�`\޻�e�������*D�8L��"1���\l��h�b���M*
V�W�Ӵd�P��:J�]#�:g�ӻA,1�Q���}�w	�@��Y۹}��޵C�^�x �F�n��j<��x��쯾��1�I������&�|֗`t=s#�ϕZú��5ᴠDK:b�z!Z�{ٮ�mh k���7٫�پ��n��W6Y>�Ә�BHE��� ��%�ֳ��7��/7��¹���P�S�N�<���%�Q�xd}�s ���ღF��u���g8���4na��M�*k#_�܎��E]w�R�?��:��er��J^�p�}ȕ�p���AY��>Eq��E���|��E l8\+ 6�ǣ1;{�,,X*���o���{՝w��B��M�X�[�~fܺ�y��:e,���"�陋(׮��Y1:F�յŅ9�W�zfh	5�o���K$��ģۺq�z��;z�.�?#
 ra���I�ܕ���9�-���m��N�G3K�m�����c1��^T�p1�$�>�]�5\���#�01d��}�N�9a�N_�=��X��3�+k���z�K��n��X�h@�3KM;wf�.M-Z��.��I�I���-�]�gNع�Ǭ�2�fi��^CH�Q�16c�%��}q:j���{������;m�ޛmp|�M�/�%� @?0	��d� ��jN�h�Z�Cub��ڴœ�X.QU���8%�
+Ѝc �n]�I'l�P���QQp�1��j:�b�'O��ꇎ���q�)��l�S�pځ7KԚ@|��ھ݆��W)�zv��Y�5�k�� nG��q9AQ�ψ��6f>�M�:<���ll�t"2q�T<RQ"���EVر��1�9|dP���J���ۧ�l���g~~W�ī�}�l��M:,fB/К��+�r:�LZP&]3�I��U� ��?]G���x;tw]��λ����ٳۮ��Zۼy�M]>k/�p�^:�����ؐr��aP�|!-�l�\�����m��d�C���^8��]�<kM�� ��3t�i��D�݃4��HI�:`�Ct;��S��J
�d�ձl&�q $\s~�l!���M#-R����A#�,fA�!o�?�Xl6׌�?��5L�T�@`:�� �����*ᘀ�A��u��`�(��WȌjZ>�@k�SFI�����sX�HY�.{G�t��H�p�^�6�B0��J�܋/>/cD��]��bp�]-����v��%�&@�Z]�w
���Ș�B2��	�W���K�d
�8�QYVJv�Y�]�7���ߴ뮾���#��̊(��n���Kʕ�;
��L'1�d ����ޣl'�_zm����Ԥ����4:���!*��*,ҹΡ�Q����}x?�5�1�ճ�O=�Q�����1!�gieU���.� ��)�+V��5�e�S�j��9�(�0(T8�N��ĦIs��ձ��A��p�x�� %2YK�s�6�p�%;{���Nا^u�m����f�jvvf���'G��^4��e|�jU��|S�.�1��*nW��kT+�w	��.�����3yh[.�\�3�&uq�榦���b��8��Ţ���[a`�r�M�I=�Hu{��~�Ct�� ��`�
��EZ��W�26>`��S�NY�� �<�~m���#�˿�s����`�v�Ri��N��s�/�r+�M�,F��b�._Z�R�vu 1����"�h+����#6?}��+���־߰x��ຈs��DF*�>Ur"�C�e
��u�u�}�5֋g��c�H*m`�jфC���07���X��֧��
�K>'+��e�)!*���=�<�:�Qt7��wh�~0��p"J����{v��%�x��e�He��	GE0��z��e��@q�adخ��j����Lr<ڸ �i�d
g��k���%,�J�m�=$,)��^.�b��Z���5���&<��"2����H$D:L�ӂ�K��zH�e�)��g��a��$�ba��d�@�y�V�c9�������Ҫ
��p�n������~�}hؘ0oBU�E�pld>�.G3y*C����Ȭr��D��a6u��Z��b��#G���%����u˄m��v�&>C�Y�L.-�*R�!R9t��l�ν�er��S�����[]Z]�:�V6��{h�gf�Dʊy�X���|{&6�Y�ӶS�O8���;�N&-��pIP&]8|���i��X����\>�{�rH�]�������/_��	�!�@���"/$+S%p��_�J����J�qrh�ԗ+�hS*x����l�g�ѳ�E5�
��%&y2�3�'��@�bw�N�;<�.R)!ew�૥�(f�x�?���d����"Uw��ͶqӤUj-���~;u悈����Q������+;��
qAQV�;���ȟ�$Źo���]������R��������������P�~�fY��HA� z���{��~���;�����m�H�ګ�S�?MG���!*�$=�\2�A鴾��6,(�b3����X8�Gy���A������|%�f�Gyfʩ�TV��Z+s��%y�=�����bg�9:���5����*���MLl�]����"�&�5�%�6�Q��>�4�K1�����뮱׽�M�ǹ8W�Z�`�Ƞ
�h�Twwȅ3>W�z@�Lv��������1c&���u���ǵ��h���OY��HxUhBj!W��ek�*�dwZ�:
���q=�*4{��koj�T�j��IN!����c���b&!��M�Z�J���T���pF�
�T��d�>}���?��_��W�����p�Z|���K�^�F!�� �-w���<��� ].�?��t�J��7���,����s�8w�je5< �X�����i��"%~�"�62��v��
�,�)Z/��F_TH6턜ÃqD�ъE�uH���t
_L��@�s�;Ӷ�K���[��J�+�-��@����#�vM�H���,�,�x�+�����DȬ|H6�����{H萈GĿ���6624��̈́�/��(h�!�q�{B�K�y� �;���A��h�k@�
${}�Hܹ́wt0��r�q˻t��z������D0��p�)#6�Źy��|pH���rpb�U���=(v�{|a���iK��x
6��M��5�aLg<�i�*͖�pn�EHl��}����Ѱ��î͆�S:7~=������	�w`�=��Gmai�Ri�®�i+���f�%�A�{&����|�v�g++VZ�X��yä�ض[c�S/�TNf�
e�e��Z׊ټmE�n~�W�2�IFhgN��TD��s2����5���{����&m����/u���݁2�C�B;�Y3t�/璄t�? Q�H�ϡ��X(�:��ٸ�4�be�A�\��c?`;��&�/�ȃ��R��H��9K+e�N�q�X<��"�n��T���t�^��d\F��ٛo����O(4�����w���<R�Y�#c�6:��J��={䈝=wɉ���c(x������A��x:k�+-�X"�c�h�e�F�^w���?��M�ڇ>�c��c�E&��e?X)e�x��	��88L4Jo��-R�}�ko���ߴZ��Ҥm�ܦ�D��Ƶ���?����2_^��HhX��|���ѹP��cU�]���c�����������`�:�oE    IDAT�mێ-V(��������td�Ui��.�8�7
J5g��J&���XH�l��-v�UW+Q�ĉË�(Au;	�ć�t�tB�$D�qۭ��w���v���ͭ"{��Nb�,�so�Ã<'�w�6�w���ذ��ZyI.�,Rx�^�]�'�¹�@JF#ڛe�q��9hp,#���k^��A�D��N,.D��V���"���b�o�
*T�Ǝ^�5�A�<�B��8,�
�'�L_�������#���-��|��Z�?�2TM<���_kŲc�%�Y4�?�`/-Y�	,��ܼ�NH��nǒ��4�"����*�l�tȕyk׫���p��b��F-?0b�C�60��,��D:o�H��p��j$�ݎ� �����i��9�x#���i!+�;����o�m���qay?�Eɭ�;���� ��̢����N��f�\T6�1i�����R˿�rVr)[2p+��Y�*6�[-˥�Z��=��	�%�A� �S2�>#���4[����H��QwX�AT=�G�-I(�WJ�N�+h��~:�W�U�
�~D�lNh�%'=����=W�ѡam��l��ݲ�.�/d��{���صS���&��J�˫����f[�T�"ON@7Aqkm.lV�{���7�%%����؈��]�������ߵ�>��u#8�bw^�D�g�B���1Kg�i3֚u.)�vĚ�����֪5�׎�P~Њ�A�6:v����.���A�����# N��U�R!���
;����n�i/�6��X�L�t�rż�����}�'2("r����}]�RϹ�y��KU[Z��b���	kы��a��a�!r���`s��?䩤SYߤ���P	a�а4<̂<���k��r`�h�|�FǆU�>���v��w�G��_��g��?��g �H�$�_!�\o
q�@���|sM}F>WRj��}���;mnvZ&i'N��-m/��}ێ�6��c�mG_<f'N��r��9;"74:�ò\�o%f�j�R��[��i����
�H�moz�쳟�O�[���Q{��oKqDSQ����-��U$��I���U#	rl��������y�ժs��E�vႫ˔�pT�*�n���6���������`�w�c-�2//H֏~֯3
I�M1?��r��7��;m���ZO�{����ʾ��SRt��h%��]_PlA���$sGw�!�m��r�=���v��A��a+��I��$eh
Ǿ���@���ko{�;U��tv��KQ��&���T�!ۏ�OJ���f�`�q.����x���4�B�!�Ie|Ͻ �w"/��bO�;�	�@�"����i_���^�G���"���Y��(O ���Ul��ذ
�R��(� c���s���H��f���,mO��T�ԯ}��Ͼ"
���˃�����;��V,�!�^+TΜ�����K�Ȧ�&s�\p���\�'�Z�o7JV)�X��Au��\aP9�)��ɢ4ku#�Le��^���v�D	B�Đ�ߕ�8���\:c� ��MP$ڀ
A	���-�E�T�vmY�Q�&�$�!閤ϠP�h�&w�́�B��QK<�_���ɟ�����euR�/��]��� {�|֕"�AbeL��N�BE����~W�ӵbqH*]kl:ݸ�=D��fV�$�q(1����̊��B��<�.+�{��[n!�@��f2J��{�n*�?k���.t�X��US*�����ط�ܹ3
�z�;�!"�W��Um�D�������ƹm�v]V�5J.�t�tA�� �^f_A*%���&S��C��W_e�~���3�[��b�cE��J��7lx�`��`Q��t�[��.� �?
f�};}��6�YiX����U�ܰ�6�L��̒-�,�h��$���Qln�v���ַ
U��7�A��7o�^��B������g�}f�i��������~ɚ8Ц���~�k�ݞ?zL�
(��JY� O�B��}�R��S�J��B�v�lpnZ圦iQbv�F�s�B���+�S�u;*�_�(د�0��F�����O���عMy6��+�l�_|���Ak��V�5���	ֱ��Z4.~x$�Ik��uh�ZJ@Fe7]���-wk��x���3R���+R�Tj5�/)�k��-,a;А�[�V<�<r;��L�s��IQ$?\z�J\BG�?�,�|������366����۷��-�U+"�W�U�4��.^�Rv�ׅ"��>�v�;�&��t��P���O������L���˗mv�LٓT<i��6�qE���'0b���Pю 1�ʋ��^?�L���ש���__��u�LN��w�!O�-�7Yq���,�ʗ��e����e���ܴ[ Niy��{3�K$[�,����)�~�����g�tK�x#~*D����TL�5łT8i�v����{�ŕ��Do9f��&*;G�h�z塔R��3�n5md�h�F���Ezuk�V�\Z�V}EH~"�rT��i�b�ګ�$Ј��}Ū�E�� ����Ѭ0���MV @��<����웰���ͱK�̐�5��Ӷ~�.2��G�K�^����4����ԯ}�_�2
���~~�k;7��3+�-�°��[(u��9����N���}m�T�n�E��0%���(�m�� w1�l���^ި5::�52�#b�a��qJ���ZP�tt s�I�]����@�ArF`M�>	X͒E��0��6��,Y��*I5�Y>����aRD8Vu�w�z��mF�-:d/H�x.���q�5�⹨bR;	�3(T����C��+����__c3U�ļ����1�^x�	s0�0��"2�0��bS���X>��J�"�*�On`�
�#z(�]uNh�#��=ldoz�딟A��_��6\�׾�ڐ�X�}�Y�����o���N+��Mw���|���ӧ���9u8�>V�V׸��WW�	P^�\��H���ܨ��9��G��d=�wk劽�-?d�~�������o��ִD�g�n�R��e�1۰iĲ��u���-!R��ҹ߼/�A(>#pu�I�F;�8������m|h�熬�R�g.�O %SUs����1��x�����zR��ؐ����[��&;��V*�J��O�>���T(]/b��������8~���%݆�X��J��B�c�����k)��B��s4~�J�TZOA���*Co�+��F���O��L6e�B^s|�ś6M��>����}���~�Ξ:mš!�5�*8���N)���()��Lc���u94�,�nw��k�R`gOq2u��҇�\���2�\Z.+C�Y�| ����ݐL꺈[ҫj�,�ˉ����=�R^V�鶔�����lrb�~�w~ێ�Ȩ��m[�Z�	q\XZ��G���ť��믵����>p�Z?����9��>!,]��]Z+T�h��g-�8�%L�#&!%,N�B��r�B�{�҄|��ꗓqף-�����-v�m��-7�(U�"2I;x����G�����΄v�3�sm�� ��GB�gH^6��"����)?�v���t�h$5��Uи*/�u�Y��B�]��gK�-;qf���QK&��F���*���d#�z�FD!����>�^^��O���Y�ڲE��k�� _$�˔�.7p񸖨��#���U�,4" 5����μ6���%�(��v�����蘭V�S�b�n�8hok7mb������*
���u[�7~�_�2F?��Ls��]�}�б��#��Flz�f��%�i�U��^�p�����1��
���B��1���Ƹ��w`M��E���q�*�@Aj �Jx6�cw������tB7in~�gg�[�+$�ҁp�1Ìźf�"Xw,��]�u>�W�%��w����$,�l��h���b�<�$�w�I9[Z)��'���� 7���k{�.BQt�٥R#DHLh���J\&a�i�Ҫx�k�w+ Z"���g&)X2 ��5�ǫ��/Ef\��ǁ�EN����lhxT)��^�
������Wh��NᏇ-���{��^�t�}�+_�t�Ͻ��eB������I�e��nt|��~��l�_�+;mwwՕ%�8�g^��UWy O˿��8���M����\�	��?�cV�U����RY�X�b�i�~��'�mh4g�<�ߖ5���d���EvĻ"X_GZ��)��o���~5V[*V&ǶZ"�s'�[y�$���Y\̋�\*gW�ޥ���/���H��¬��ۑ��ZeuU�x?����?�Aڂt�~H8p�N�8k��]Pq*p�<��+��c=�����AW�ӉP�6x������'v�"@T�\(���$�""�e�!)b1�����?��_���&�������s�-��Y�ٷ�JM<��hV�狍;n�DF��o������`Ċ��]��,��P�`AyD!���"�$�0{��R�᪥��f�#���gA�h��y��d�B�Z� ��?|�\.e[7�ڞ����2̤�6>>&c���ޭb�ೇ�~�]w�^{���=hC�BS�c�3��O��R	ϳ*�υ�R�i)PhYA��J�����pT#�o�׊FP�u����I���'͆����~�r����~�v�-�ڮ];�8XЁ����w�5*�A��Q���F��F�42���d6o7�|��j�������=�u���ƻ��Q ���Ka$���M7\o�y���Rn۱��6�صHf�ZVT(.�!́q&?��M1�4c����,L[*�ҴfgO��3/�5W�O��&�A4nQ�U5ZgBS�rr�P�2k��'
k�b�9�t�ɹ�ũT8��ⓤ�r��6�q�-,�j�P!��շ��P�����HT�7(T�����������W��g��ϭ.�������/^�Nzr6? y�ԥ�xq�ju/"�P^�y:.� �1,c*��\� A�xB�i��J���������b��9���.mM��=�]Q��*}z4b���;��	�4� g�Y��ױt���[;떼Tb��eS�{�ps@��7�ƾ@lJ���(2�L�X�ʆ�44:&8�¥)۷�;q*�$|�MǨCA;?eAe�Q}���8&�̷���(N��SԦ��h��!H�Q�7��շF	�ND��Wm`�m��J�2��Ώ�O���%�L�諃��g���W��d|-��w�[��g*����O#����Ry�n�kqa�2yOÆ����җ���؄��䋊�����-V�4�$-�t){|ӥP�H�4�H%<�C&IJ#��=�y��|��O��;s�E�\���[2�������L�a-܏c���N�t��f,���_5,��VY�Ym�b����'�{�bO]0����3�j�t�&7M(�l�����"S�u��{�C:Զl����?c?��#���+�Ҫ=���ꬉN����Z��RE�)�D��u�~a�)a!��ZAbv8Tg�i�Wڠ�[���;���/���.�H�J��m��JA$T8U۶o�O|�W�e?�����'��rm������\r�!EILO��5�ɠ���ճ$\"d%����Q1az0cO�ͬ-���_i?�����B�y2����^]��,W,����Vr	=mBɵ�Mc֬���+�Rʆiԫ�m�6�!d��uhd�n��:{���w߫�"��D�E�}�I;��Y��C���ȹp�9,f*n/�Lfn�S�>,F����P	����%,bBt!��P	��^��ɍ���[�[o��v��i�[){�'���7*T� �iu�J�G/R��ׁBgr6<:b����򑦧gE��4(�p��ZV��-?���������uo�W�x�*TJծ?;k����MZ+:h�xN�:�ib>�L1"6ۃ�`&�8s��Z�N�x��N�`o	]�[G�8H0c8� E��)^P��ԇ^(�.u��ٍzH�gn�}(2 ��Ę��y�޽62�Ag4��l�я���P�<9f/}�^:��5)�R �QKZ��5���o�����WD�2?�/,G��}����6�z ?=6��pa�ʥ�K��0�p��Ek���T��/�<6{1�{~`� ���x�f��4Dl"�<��\fR�(����Q���Z��l��%[^�wc� �Ü?}����������KmT1��G��al$8��l�U2�p|�L2�f̄_�
dZ65ȴ��!�l�Μ��_|��I���C�{��� ����	VP��C0�|�Q�|��I��~m3V�o@U�$����$�txD��rG���� ��#�Ctȃ#����#q�DB넕�dUFy� D0�X����-����}633c_�ۿWe`h�>�������>g�l��Q5��ղ�r��]w�)�O��*p6NLh��ݯtn���ВH��@�\	]g����k���I��?�!�6:������-��Y:O�ж�P��7Z,Ł�REJ��%��aK���9�	��2@�X��:EpªK+-T��P�N�kG7Y6���/Zm�&"��%���٦���g�a�׬Z+�ޫwۙ3'ģغu������=�S?�^A��]>����Gmnn�N�8m�/OY��[Z]u�Ȉ��:��Q〰���9o���@6����5�d`�*a7.�F�'�s�k�?<���hz��c�4juk?��_�[o�Ŏz�>��۾}�솛o�Z�'�+��"O*h)=�qwF!d<�q�X��=�Z�>����$�oY�;I;�p�(��c;�3F�[3��G��f��P�**�o���2VWe��J���,Wd���&h]�o��=?�}�~�����̩x����o�=����o=��]_�����v�د��ׯ�+G�����p�6��Ԙ',T�u���֯��P��G=P��t�M2�C}�g�U�������/|���?���$őHJ�BtW�[��:�����B	���!�6
�B��%I��N�Zq@����N�=��F���{�}��V�v��M-t���-�<�功u��k�
Iq��`>'�~i�����V���p�Y��4�5�V��U�k�ǊkME�C��c/�h`J��`4���p�\`��C�e�V�m� O��h�=��*P�n�`�<m/�8�P�d6��/e��WO|��}�O^{�������������b�o�97���*[�W�Zo����/Vlff�VWj>�Q�bš<y��������U����![��P	T8"2��L�kw��Z�⮚\��Xal��IG*	��o��
-��t�f�g4gdQ�|��G�Qկ~�a�d��J.�XK�
��\�R3y�(�{`�[@�@R���A�#�h���GF&��B�1J�蹞�*�OίAx^��i� l̌(���A�5�*�@d,�HUy_V��ս�o��o��:�Ɉ�������Ç���mۺ�햍oج���CG�����ֽ+�B�C��B���܌�!����g�g��\DV�??��Ϻ=?�M��p{���/���̟��T�nhu銻*3�+�J`'�.K&�u@��	��Rph������f�߿a�?��e�	���t-;�M[�-�9iX�UV'�g	����:� �T���(&��N�c�^�*+u+ϗ��P�L,oÅa+-Vm~j��-�-�\6g�ZM�����eKŢ66:��diaF��(8G�.�Ͻ����s�L�mO=���(~�,-�� ��>��
�wDp��6ʰ�]�a���</:�l�^XԄ���$�K
|O�Fl��*�NH��r3 p�
U��䐿���l���ZW��cG�<o{�^��
o�sQ*⯏��QL����p@��WA�E��E~mTF~H�BJx&C�+й�N;��ȓ����'�B�ј:Y�s����bV���Ө���k[!KZ�ҩ��,/H�i�ƥ<��'� ��*qƩ�}�Ix��s@g�ģ�+-yxx���/�R���s��ɌD4]��p�B���n�^j�& ��o��H���џ?ڠ�W2{�?�����Ex���\k{�챭�[�n������w�/��W���#ڋ��    IDAT�Q�FY����8~��"��1�qL�sLf4J��պM^A���*�.L1]ѳ4�T��2���.[)7���E�Z�Z32 ?
���|M0NG?*�[mKG��`�\^�l�8n�-��|Ϊ�y�P"��EF�}5� �4�<� �1�c�f.6��"�6�s2�x`2�'�ʬ_)��	D#V��e��L%,�##*g�|ڲ��XO� �?�tl��Mv�'��/�P�rRi��uy�D�w�g?��WD����|�w�w�7�Vړ�̠�j][*�mf�d�3�67�,EĲRW
.n�T|��#�˚��p�IBc����n��I�H��w�T�ghX㛈�]蚂�������q#���%đa'��p�����V+�z}*^\@�*�Z�Z͚� ��(-X���Y6@���Q��ۏ�俀�q��)��Pl:�m43g'	X�*���X�ڥ�sh\*�5�t']т�ڠ8�I�� GE�!�V�!�9[I��j�{�A���7����_�#�������:b��/�!?>��jt��m޲�z����A����O�a&�PQ�7���=g�Gq����{�{�����_�����
������O���¥i�w�v����?.��7��u"T~��_����ܲ�9d��Ѷ;�s�U��TVl�`h�b�'	 Tv`�����,�V���>�ÊJ����'���d�Xˢ�O�-?��P�i��R�px2�b#�@Fe�;a֢PE��f���ݾ��M���iFl��J-�F���uv��ekW[���ځ��a6��8�594�Qyf���*C3�b1/�<�RܛJ��S,U�#����� }t����	E�����G��	$�M"�s9mb*!2�2�9x�u�ayd�4@���v�c_!P��S8�u�.���xp �b��1�?	
��
��
�1
-�2PH��MU����_rL/�$����q��z�8�$w�e�#��p���ƍ�zvc�K³A���aߜ�e M�Uk�];&miq��f��������֭�%Ӿ��{�����铧���i�J'���<|䈊S�s��8#V)W�,�s����$%Q�+��AF_A�y������B��c�O@�u	E4�~I����c�Ȍ`�V� ���$,�̯�m۲U"��^:n���$Ő_�/iu�o��������!
����q5����a�~�["j8�4��3i���N{�[�j�+%�0�b���Y+2l�X�_�x�P�S�� ;��b0@� *@տVW�o�UT�MSW�P?��V�g֌�u�4����'��R|$�U�[�qQK<������\���_��#��}������f�*�sMq�"ֶ�Ѽ~v��<sҺXd��0S�|�Ɓ���_~����
@Tί�U��7?��󟪷����e�6�\��f��;u����]���J02Z��#�
*���Nb���P�x\8�j�C�4Tʉ't�ʟ��.nb0R����qH8�&�tr+E5ĜOr���Q9�fب�\��	�W #U���q�p8�
;I�Ga /F9ˊC�Gu���2uj�I�R���BYg�%B��w6�]�,�9A6l�� ��zl�\�L��$눽�}�,����4��u6n�l�|N3�0��8���Q���R��?��?��G�����M�	}282B>�$9�B��7��u�x��o�b��=�)0?���̼��i����O��G����׿V���G��V�R�5��}�n[Z,i�d���X��W�?�R�@�d�q{��iS�ҟ��U)F=K�6�u�
���b���HKǁz����D�~���*����f�
E��~p��.�t��*-+ϖ��P�N�gùQ�%
v��%+-�E�Sw�wg�l&-#�\0�i��v��9�[�,hM��A��K�t��	�K�R�}ٴqRrf$��|�m���xM�y��*A@�EH� U�\x��U�� ����#��"����s�n�$�;���I�al��$��;����:�l4�y��x٘e��Є���R|�m������xr�#�:��{H,��P��òi�.\�g�4 
7��ϯηz6y�2�ž�KA� �C{=K��E8aK$�˶c�F٭�MO)DjJ�c36:>.)��౨B2�A#�Ep���S���J�r^	�
S%#+S\�1��3�(�Zw�c�c^�Î�f�z�ȯ���"���X7���X�{�	,�6h�v��F�A`cW�R��Ƞqm4dT	�?�H[~p�Z��+vI�Z���K�+2=M����I\?�� RC�@YU�E���%<�� ��H�n��{���f���]�_��=���֊�Z��>v!�V��^�i��r�	����N[�=�B�1�W��tJ)��x<ݝj-ٷײ^�b����
(P�`�UQ2��b�s��J�j�e�-?8f�*����x����8��cdt�
����< ��:61V�������ܛB��H��5�~�?�ӟ{E *X�'҅w~{�s�Ui�6o�n�Dޚ=zy�bS�Z\tq|�P�0�Ġ���L����`E���h8!3`�á��I���X��5SU)��F��� ����kS���R��S���tt���/�M�p�3��`����/Y���9ߟ�x���)�2}GTdO���?���XV��҉� ��aj*����K�0�f|$��ЫA~x�!aT��Yѯ;*�[8��0hU���EZC�g]����_��?�����86z����"xqQ~�^w�=������>��wܗ�׵^�������i�u-n��V�{�]�c�^����d��(�-�;t���|����S�|ГZ���DڋB>�ɴ]۹{�-.����%BE�� �%������G>������ǬM(c�m�Ѵm�1fc��lyeƲ���si��U ��BTʥ�U*e%�B�� �*V��k6�~�c�n��+5k,5le�l�z�3C6>��Ξ<g�S��*�>�\�'�c�����fy���0�Wh���Yn�]�-�-���C�3�y�7�	d�/����)�����3�Se��f���J��B�tt2�':r
g^%(��8c#A�~xHi"��2:�5X�Pm�i����{�À��VߊC�*P����Q���c0��p%�*�P}?�I	�(*���e�+#Ş�u�R��$�Ҷ��x��"-��ED���&E9�i����/	T�i�7+T�b��?N�n�|��U��T�.�8.����ٱu�Ml�$#E�+�Ό�@W��ʸ2�ZEqJ���hD��b�'��}S�3�4�:�V�4��H�@/TPeʢ�ɸ>��B�.�wFj�.zp�{�탵Ĝ��5�S����=��r5�Y� ����[�1�R�UB�����pl�:�L!���N�Jَ#BPT���nػ���V��mz��B��/Z�?l�~Jd�>5��p΀źcd���u� Q� ��Kq2��^���8�����Ӗ���QZ�|6a�Hώ9�U�%�@�\q��ɬ��MK��������b��m�5�ݨ�Ղ�Y(�l8��x�K�:��
��C��S�����;M���[&ھt������W�{�-;���g?�e9*��~"Ϸ�>��r=�ad����*T`AS���.�PA���!<@����"��u���/
	eϸ����q�{'�2�e�V�X`��"�3I��[�z�XĪ�����y�4�}m������^fL�uU����"%��۰h�1p��}�Z��$)']7�:6�Z���y*2}=
}��b����k���>Ur[��e��	���1�ps/S)m�
�R�&;p�R�;z��*(��ldQ��~��O}J7sa�<,d�!���:{���h��L���E;|�y]�zS�0�R6�s�y�?�0�S�X���9��,K����?JO�E�B�S,�!N7�hc���H�91�I�5��`�ݴi� !*t�w��u�I��Dc���u�����}�;߱��;����-��D�&���H�
�q[Z����`�n��z��l�����蜃^[�]���$��s�j�ڵ�u�mk�[V[jZ��^+b;6ﲓ/����Ӗ���ɣ������'�S�٩˺�:r��ޑ��p��`��m>-�2�Dz�5g��F��C�۵\:�#Qe�D�.àH>��̠VK�+�:�Iee��z��R(�{�@�!k�<X���� 84���	o�-��N��~�
㲩�5a�� SRv�Q��
A�����
�)f��(D��ϕNk	5!jxn�.WZ��r���'� �p����RA�r��=��b}b�1 f���T?t߫ˋ֬Y�e�*ݠ�	@����<$mh`БF�ф呝f��BM���`>w]�����~�jy�G���wA2��JF�h��Q�gfR����|)�د����CK�K���UF�ڂ�g��؉�coT�����T�%)���{TE2%'tk7�	Z<%/
UT^�6#.�7
���Ta�4ɣ�I��� ���]����񎷉�sqv�.̶���Y�7dM��4��W	��
dF�15Ɍ�U��k�����s8l*�G^ĉh͈'��B�z�U�'z�8uά�j�#�Coy�����M]�� �VKZ4;`�lQE���[-�-Z��T�FC��L.��^ϼ"+R�u��$l�H*5"������R�<��w�
�Z�r��k7��o|�'���w�Z�g�� ������_�sf�����G�܈���J���՚-.�ly��nU����`�⇆sI�u�͔Etᘌ��&�͓�}NHN!<)I4�΂���/f~�7� �}ѳ@K�+������Q�9#�~Ϛ��~�P+���jV+/Z��"��>ԉX��̃�D~L+8(&<��Ϥ���_r� :J�)\"��g��� �u^��5�.�#6#d��{3}Y�&�@^Kg��86d����M�kU'����l(l$�<�m߹�~��[Hئ-[�	�#����w�c۷�?����c/�~�e�*Uu��f��QKQ"��g���!n񺼟������O��]�T���cӴ9@�Z8�	����Ai�?�3����蠋#�p�^q�p�a^[�N�#�	�;L��;f=���U�4h#y+��l`(i��%�=��5����FU����씔8-п(v�iK�S<�#ĸ����ƭ�ڴ~#j�~�g�����KG����b�g�#?8*gsI�W+�U�4�<��?
�L�@�#UW��a����'��&/��F��)aQ'�K�U`!�cH�/He�{)�a2c��l6���}���"ۨ�ř���u ��q�x;�*mM!3C����F�C��ST��!�} Gd~`�b���=�t� ��Eb��d��oI��GE6^�^<h��� VY;�Ln���p1(
A�Z-8wA~W �>B��uV�@�T�1l	2�$ƃ\��m��@9@�A@@��c�.C��=��TRJ"�����;���a��s�ZMg�B��QhSW��u#΍c�TJv�"%S��+4z�Z�?�3�� ��p$f�thO�����l��H;P_�^H~s�U	{�JSc
��ٖGH�(�c�ٓ�D�Mڸ��8�g�C����(��x��y	��RL$!��7	/�B!8��ݯ�����Rȹ�;7ݴR+c�ޠ5�nE���"gYO/�Q��a� D�j���n�%8!}�����'��Z����a| ms�NX�[���mb(c�wN�C�g���w�?���X]m�d:�k��rpuR�t���l��vK�mn���Od��SNéCL��5���{�2��З�I(c�6m�}��kgϟ�N�	��8��ū'����FJ�3�ſ(�rt��!��=����m��-�MZ,Y�N$neH��e�pqFɢ-X�}�9���A�69 ��r<�6�P!!���R��� F�Ε���8�BZ0ـ����@�V�lvzJ�OWnB��!w�;T���O�t�*R��Q�t<��ߨ�3���!c�!u��S!����Q[�qKR�*re`V A�t�9b��� ꜃:p�,����acA�A63s]�hT��gDt�������I\�-�0�^nr508��=���f+�U�m5E���>�>ٖ�3��_��Y��$���H�QO�x��\%ϻ,u�̚3��'T:�!u\7�Zf�@���yJ-�$�"HZ�>���_�
(O���tN܌�@�A�8����}�����>��
�~�a��8�������V,BW�cW��a�^�W�n����[��lj���1[(j��.L X�յ�Œ%-i�Ū%��v�67�d7^{��<zܦ/Ϲ*$��sE��"(�p���)qO��<C61��7�c](�-�K��2x-�dC���1�9x��@��Ty������2d��lanNk������π�K�PFH�ʈri.���w��.����E#�E@��{����k}�" t.P��uB
C�#������]�Y�ʀ	dGz݀{�dx�^WWhD4T��𱮸�H��9��9(���l3��z�U�.M����EM�s8�u�J�FrHZ#�j��\�)�JyfX6�C6���E=w�B�,R�P�4ߟ�����g��p�8������i
�}��Jc��'�_���	���d��$[��|$�gFf���<��B-��!z������#�!/�]]�aKAzYǄ��
�0�r$==j}�A���p�e>%Ү{0�Y�̪$h<��o�^D!��}���η�M����Kva�i�nњ6lM�@Jd��>�0uΘԖ��g���G~N��~�Lx��aZг�B�"�U[�?k���M{�Zu�E�U�n�.�j�v�뮻�w����z�*���'���D[k�^"���-;l��k-��F�o˕�5:}�˰)�{ݺm������}�t�N�E;66ZG����@�e_�D���(|������+�Pya�2�̃O?��ǫ��(dZ�e�ً	Q��[�ٹU��ڌ�ܴK�@�"E�Z_ꈵB%�v�
s�`^L7�. M�&x�-��G �`6��Y*��hZ2gc�ݲ��y�|���`ไ)�H+��P����-i���ي���kU��ƣ@O�H�6oQ���²���Iu��xA�b�M�Vw�,�K�/0��t�g�!��kf���<��h�eO��4��>:��7��b�������U�aK�͙�rju�����i���[�xX^/?�I,��������� �?��?�@3q�"d��� ��b�u��DN�%ח��k���T�c<�Q�����&si���E��	R �,家N���D����	%�d�N@�˹��oG�|����ۏ�؏����Ǟ�/-���0����F-��xW�V�����-��o~����;����W,�M��Ϛ�Z@d�QTE��j���=�T��<W�x?c�R��c��x�=x��g������6�LCAY�G�Q��u�3�$�С�J�!.�b�AѨ�p�4�%�[u�� i=�t��Zv��I}_D~�`;���hp~f�ffU�_�����N�7�$h@͎�:m/]�{c���*��);rL��y�!a�έ��H�)�@�`��g�qi�dFExr��-���x_��w�Q�$���U��@�����1�U��a�B�t�:	��Y#�`�Ğ%.HB$�ɖI
=6��#��w��ѷ;{���6��{t��)���v^
9;s�=�}ڋ0�� c����pI1(��;�+ph�����C����X"���bڻXw�#�G�}�Yq /e��&�.��x�*h
���
w�HT�
�-����wo���p����s�.\c���j������h�T��l=��h�<�����P
O9):��Tu8*�7 z�S� ñ������{�!d���]�oY��S���g�d��W,��Z\�0�P�[i��X��@TجR�`�pBO�m��v��g,�^����}���#�m����f�ԙ3������Vkvmn�au���s�v�7+nۮ�ή��U�����e+U��r��E��2E�<>h�9H�,�    IDAT%�R^r����޳᡼8��?���PeӺ��~��U���7���忾b
�����̑�~�҈�fa�G3BT�KM*ӳe���Z����<s��)2���4�Y*
^�$�nd&�A0! �t7��Er$$����Q�C��Af��x4h�Օe[��U��S�h���PȻA̹6�NK��*�ʒ�V�׮haŌθ�`ūw�V�������I�lMr�M7jSǬ
I(�Q����v��a���K��7 )˩�l�!�f�II�)H��x6��.@��	|0�>yۮ��λ~�����0F��p��29?����=7(j��7�ٶn#+gU������/h#ڹk���'� �:;�Yϐ0%:#�pH�2ڤ(PB��6����]�(��9_A��̕�s��[
1)/��u��߬t֠2	¹T ����%�nYq@���/��\��l�H���q%�~��_�6F���ٵw�2Y�c�"��%S��^�w�x)�tF=��Kj��RDc�N�-��N�QkX:���������)��]���v�k�{����������3������J��
B�c����0�rN�����8��B1� 3��i�+��\�9��4�|��w�[�ے��y��}�s����9,��������	����C��?�3��oî��{��֢���WV��կ���D���5[��&˗}�RŢ�X΃�PȆ���Q�].{��&�e�m�ꁷE���32�B�OCwB9���Zs������R>؏>�	�!s����B�C��9�'�Y,�*�ZH�G��E?̓$Ύ&��;�Goj(���qEVLn�h���v��]���|��Oأ�~K?YADQ�Pr�{ _���=mw�y���k~@E7�Ŷ����g��N�9#�,�4�E���h���fw��*����Zb<�S.��[u����F�{��;N�\/���M��Z��6�APf���a����M��i�mب덏L�8h�|޾��3��3�aa�.���4*�\>�0Am3"~q���Q�d2ڵ;���}�ۭR��Ź;7S��f�j�ջI���H���Q��0�e�-�r�UJ+�I�觥�����\ڬS��K'��ѧ̖/��H�>�S?j[&�K���64�S���۷��?}�.ϭ�����j�mMԨ��-���ul�-���o�v[,�mayբ��~��l�c[7�X1���Ae�ź6P�ؑC߳OS��>O��V/�(��'��/}�S�D��<s���-ף�P��Q)�����4W��e:��{H���^-ɥYP�*�F�VV��s��8/Y0s���� W�������3Vit�� �&oq�"�B��jW���gW!��,/�<	�x$ w��MGC'�$9�'��w%�][�F��R$a��E���j�N�ת�0=��0U7p�޽{�G~��R��`!�'��%��?��*����XYXX�Bc�6=8$]n�9tU�k��fYI�|*H������CG��sg/�DV�7��-��w����\�T�<Ԑg���00hã�:�J�����~Pt �!S�ȴ�k�Ԯ�Ef�Z�y3��0�aAm_�=���,~��`���{�(��;[xWΡ�s�V�	e!D��B�d���'p�y�z3���}����m@�Q!@B9��:���9o�έ���[���GϚ%#�[Uu�=g���AKo%�L�&<�*��ZaY<Ti����ښ����X��e�����iZ�1�^�(I���ŤG��Q�]�/|�N�G�D"W��`�Cg)`��&8��98=Ԫ�`��H��p[MD�. GKL&P ^��A�Eu7�L9=��,�{�p���8x��8�ԨS˪ 5-Y0�0[�����a���C�RP���Q����S���
��i�(l%�%�#ɬd;��o钅���+��_����=/vr2��tߗ$v���b��l�eŢ���Ʋ�Kq󚛄�:����w��8}�,���ZDb1	;$EO�,BI:7�N#�*�]A�t�6�1q�fq-�����+)��|�)��g@˴�8�#?�Raڴ��8f"sG�6�ԫ����)�~��bф�Aa��&*������vfj($PN{�d{���wv9�G�KAu�����y�� �_:#te�r|�ѝ1c��.q���a����%��z��[o���[F��/�M�yE�'OFUe%6n�(�)���x�1;y�<�<��$T�Q�fR:j2���c��va�wd���%"�3��n2��f�OZ�$�р�]��^�V�d,ȱ,�ɘ��#�B��bJ1���k��|)dUX������\�-h�8O=�Faē<iQ���ώ�8�#�L��p�>��@����2��,�3�ܼ�HD@A�p��	���dJ̅1����>J��ɤ�pڜ�8F�H�P z��Ѥ����#�Q�سm#�>��qT�t��+�����g��ɓ'循�oƸ	�񪬪Ác���!���<�3_&��a0A�`Ĳˮ����p���H��pq�y�n�u9TU8�P�E48*�=��r^�s���]8�Ӊ#ld�0�c}��~�/?�ֳ��B��Y�����'�O)G?*����7A8�JY>m�`��2���T��X�Ght�}]�#�#���V6�B^��r����U���	����pWK�K����`j.HdJ�"N �
,"P��@!n�g���v0Ҷ<��P�o��o�J&�r�IZ���F�$��m��s���+�"6�T@{k.FF�R��Ά�8��	�ˋ����ȱV���zx+<8r�X���2s�t\{�*�FѬ����I��G���?��h�uM�t�J|��V��"�y����%��	F�UT���1�`�7}��tG�y���2�HX ��	�ک\@	�.�͑$�iY��j�]P�Ҳd���'��%O�,�@J�A�f"K9�`\�E磬��iCj���������ĩ� �-���З�b�r,^��o|����j@��FQ�E]c5��vTֺ��E�7q��G*�ѬC��B��%-���� &J�L0�,��2����+��ft��a��e�T⡨�,5�N�e{.7'�$�T�O��Ha�^ �MHy!ׄ�<-�s�)�c���d�p�B�C��XM�}#�[-�ʃ���W���<Gd���Wp���ͯ�Νc�]TڬY
y��ATUW�f���#rKs|�A��8	���cpdX�lj��^���J	O#��BOqe�w�`"T	��*����	��|T���/�a�E$�F�Q�dN?�[Į�<���܀ӧ
�x��q<x1q<饝x��r����M��GV��F�]�%�R�0F(��z=R�J���:5y� GY�4�^Y�����N$�RM!��(�n�Sᚪ� ���<�-yF���?�sJ�#?$���g�F*N��*���9	UK�Ƃ�۬9�����;��˯�$.*�J��rsBF�����|��~�	�xX��T4�"Mf�$	/Y�D6Y
����_������#��*��|}b�/�EoCˮͪ&�pL�&�J˵��B<��5��ǲ�V�^���^� V����(���Sxh~��T�F5����5���G�5���A�:;�:��oQ��5��l���"Z	΁X,"{����Ȣ�i�M���{D@��(���<FT{l�ҽw�}�u�V)��f���_e*k��'�Y�ryD��?��j0��]{1N����E�Bow��E�f�����Q�u���B,�"��|
>'�ۉξn����p
 F�����㟏я ��=�O�S8^�qV6Pɖ(�U@�w0�H"}��[2'<�)���ݬG2�G`��=�04�-��ȭ��fX��oy�dr%������L+*j�Q��wULv� FҒ��dFx��EX�pdh2I���*2mլ�dTT$�?S��/���l2$�\2**|^4�u�	��-TD�[PH'�p�l�r�-�y=��RSY�Ɩf�t:���q����V�i̚=���C_� ���yٔK6eʤ��ګ1}�$�<~LP47"�&666��3x��p��)ؽ>,Y~	6m~]��2��1k�"l6R�:�m`�*7.R�xL����KS,�T-f8l�sG�3�'Y��r]�˄"8�0�� ԩ֜-'AJY�U��������YO���Q��r���;�����V4mY���@��*��d������fT^���z44���އs���wߒ�t<�[u��;���Lyu�%$�1�51�@��]*ёF��M��¤Xf���a6��4{%1�e<ښ�c�ǻp�kP¤��PyY�E��W9?eᦢ�CĻ�dd����p��BD�Cu�k�i�y�H���"�GsOlv�"����>$����_02< =Cw�~�͝-�hڲ�E-���

�u���cŊX�x)��[�w�A<��3r�exh,䑡���6�Q��
l�a��X��j)V�j�^�r!ݮѯh�O��vQq|�&�j9�jilč7\��K�k5S�lǞ={����{��^��}�8q2Dp�1���ob�';����sK�z� PTcl��FH���@E�P������h�l"P@��"u��@�4�jL�<k�Qgv�?���Z�@&$���-7݌��f��W���'�k�Z�ٜ$w��̣n��H��g�u�F%+�+N'��&��C~��G��{o��߇�l@:E:��i��ys��)�Q~WO7>�χށa�_�z���λ���;��o�Q���K�1%�kiFM�V�Ӧ�}E������k��p٪�p��w��_��#�E\Kw�$UP)���l3 Q���{T�	�t��X�7���@P�J�?�фiT Sr [P,�h��k-�\&+�m,�T��<�37��F�ǌR&��[�C62�J�5n���0eb���h�Ξ�DO_?JE�����`s�`��!\e�ڮZy%�,�������ũ�0a�B,�l%�Y}��(=Bt�Q�u����05F��+	��.@���)VT8�rL�t��Z�/��G�����oO���Qq��?Tz��!�V��^-�2�7Ұ��������8�X�/ ;��D��S�H	�^_�T���{P
�(�!b��Tj�@u}��`����ꐢȒ%sZ*)��B>-'��ߏP`Tnx�sR`��~��Qc  O&� Tr�0ұ riR���mv�4��ɢ��G�6��քkV����Sp����jS!O�*�6c&M�����`�+1��]�c'NI�嗭�h��Ш�-��㏊�����2���(q�Ǎ	&��V#K�O���ca�a�������¨��m�'��6Xe3���r4nz<P�ff�*�;���RZ`bv".����Z��������z��Ę�"L���)��5.rr.��8唫,~�$�
^fX4[�T�k����Z�[(P�/ H�]F���%U
��z���.T�X*XΏ��5�8~^}�e��<+�N�c�u��r�he�Z�6�*�H�#��2¬$'�^�!E��i�7�P4��!�¾�<��A�,N�����ǝ7߅��al�����X*F��Q�<"�dԺhN�j&_�h�t��IT��v��k],
�8U�)tL���}�cCV@�f��Fm��7݄��F<����<uR �W��e\s������8|��r5��n	�(�c���݉K.��u�X��+ؼ�#"!dr�e���Q�x-��\��Q:�1+`��cs��<���dS�/W���)M(	�b�&aTґ,+�^u%�Q|�����7�_v�e�6e��zO�<E��o��6���/���o��i3��1/���E�-D�KG�[f�@E�a���l��ɵ��h��N�ZD��!7��SL
��jBϠ��_��њ��~="� ��f�j��6�7����7���MsT�V��T���:�y����q��Qq�H$;M9�A{:jk���7����lƦo"���P�ʚ?{�$�on�BW�%1aO��0*���HfE��裏a��������� ���'����B08*�cִ�h��W%�M9���^2��-��g0��c��+p�w���������0����8,y@��K+�ޒ��oT�k�ؔ�]��K���%�n��2�
��3���*ye�C B}���}�l���+r:���C�BAgB(�qsq8^1��Yr�>������Ϣ�cA]��[�p�]����}���Ξ^��1��5��}��H�-p����1u�T,[�TFC�k�������0���Ɯ��ᨬC(�,,� XzJ�R岊��{�
��hT(�~�������Z_��'�ŵ�>9**������ ��	P!p �Md�=0*@%�U�t?Y�K�CF_���q'�@,8���ԭ���lيƺ:ur֕d��B8y���G%m/W��߄$��QQ݄����X݈�2(p&Wd��
/��@eth�`@R9. *\�頑�[�T��vZjˣ�TX�|&*]�tL��A�
�k,�Q_�]����d��?�'�Y�5l\V�E�ۋ�W��/��>=z��0:�{e3�6u&¡��lΟ�;n�A:^�=��D2	���dӽ�λ1s�x�]��m~_�Ä�S�q��B¨��D	�^T�h��PXj� 2�]F'%�M�\��.c�h0 7$m؜S$�����ڌ5��8-�hQNc�kGK��:�$���R*�B�)��b\�����xPmC��YؕX����M����!�g������o��Q��)2Ee�P���{�������W�x����+:Ń؜t)`q�f�@�� /U�&���L��G�l"�\��h(�ŅH0�X$�[n�K.ǋϽ��݈0͈�E��K1��^d3�����á�W�q�&uky3JL�S-��"lV�lB�F�'s���M�}��g�L���D<����|Ӎ�x������/܉ٳg᷿��8�qF�R�5u���齶�}}}�12��+^����v�ۃ�~xv�@N���~Di>��\$h����WĥQ��[�7��vH[�����3�W�w^��RCQ����n�#?�ɏ����yepkK���\�u����n�:l߾�I��g͙�_��W8x萌���}L2ߦl��Y���^�#��!�b� 7y���Y�-J���ʡȼ&q�i|�A������� ���S�8 ~�!�}��G��5��Hz����a�ڱ|�R\��J�����y){$��a�#4Z����#�����y۶n�����[0�����ME������V��Q��,fΘ���W��w�d����+y*�vb����0��>�=[̨��B]}-lL�M�$�B�Cǎ��c�0~�4���6�}�u;}q��2aY�&�ĩHe/�E�����4��� ���0�����07H2mI�D*��f�g�#0܃hpD�'6�W�6�WU�Ë�@i�dI��a)��o�F��QW��RB]��_u���R���+�nVTU���Cط� *�k�1��}���1ߒ����6--��?�����g8�dA���30u����'ItY��+<����X~6�P����$��g�\�
�i��_��G�~C�v����O�	T�%3��l������!�S��.�|�)d��q��N�zD�c6�`(e�q���� v+��-�Wƥ�$8g�\�4��M���@��S��p
�U��hlj����p,�LA���6�c�d��ʉ�BiK��Xfy#��%nh����-�"SCSȧ#H'��ˈ�aoI����&��9��r#��{1}�8����5��Uze\�hz.��&L����oc��Eg_�h�E��ї0y�8Lׂ*�]g����q	H!�qM��I��{�I����-����-���V���Ȱ�M�-����Q�w:��4zZ-c�R��,�\���$��t�� M˼.C��M{�/*�̚5�;5����EsJ�(ŶQ�O�d;��	�zQ�k�Bm�)/�zM���ٿ�*IU-���C�v���/�ĒF�|0���$�V��~�ʕW�"�9�    IDATk���o���|�"�5JL��#�O��0���.7O�q����p�˫9t�K��)�ZQ*葊&�M�Q�Eo� z���|�
�y�=�ŵ�M��bD2�Bͨ�&�ʱ�����MO��t�h�J�}z䊌>W �_r}�$�W�Ewwj����К��6��$��jp�7����ÿ���W ��݂�n�k�>����$��c���zL�0Q?o�gN�������`s��ǧ���'Oɉ��r˽�H�5�)�"dT6��r\ J4F�B�r!��3L*
�(vF�KX�2���.�Sґn��6�w�=����6�'��==�V�E��V��O�˦��Ԉ-[?���#c�(�i�k��:7��=+����Lk.�"
�(G�b��I�"��P����T:�,�6m���ozo:;��8���#G����[Y�+V����{�g��n�C;w���r]�RDiq�P�$��_D[S#����x��cۖͨ��@���-�"�6R�FCp��\��zQ]߀��N�}�x9D-X��n� =�x��'���xe�+p�X�l���SƵ��q+�w./l0�ݙ3gK��P ��m���ª�k��7q����i�ؗќ�1�E�t8&,�Tt�r͐ɴZC؍FC9��+.Y"]?�s���0�/JԨd�����h�?��HPH��V���H�I,���Ar��u��x��W�LN��5�5�bbk#Z[���c�M7c�vlٲ�o�P��(ȡ�섫�𡿿�^z�ܳ_|	�۴�o݉��� �ӣ}�l�]|	z��(�V�[�PqK"h��5�T�ʚw��}��������)ޟ��'����BL����d�w��b��"˄ͼN�J�@ �q�̖�����y�Fp��A�w��˪G1�+��q���x��k4��V)�Lc\0��z�ܹ{�@IgAQO�	�X�0`������V�K����W�C�˦��B!�"��5C�t2HO��0���1֥� �,G?�
��W��bT�ҡA׏��A��������y^�[�-Q:�P$_U5�,_��|�=���o`�}��O1w�A��.[�W]�C=x��������QWW���
:<�����ٍ6ax$,��[>���(�a���7��/���$�:�H��K,f����e:C>��A�&�X�#��]^�
w�bE��3����ɋ�ʝ��)5z�x�,4�g�5��4�f������E �7j�c��d�� ������)/�b5��Pt� 0@Ͽ8�0�S.Ga�]l�(V�U�.�_��#r�ܸ�=ؿ�\
n����p:	�'�W��hh@�X2"�����(�O�"��"�ʩV�h5�5
��m<n��.�d�'�w���_��@4,'a6�a #E���~� 0=��b�e�G�nh-�������`*-#�f�76`t4 �M^���j0�n�M��
,]����By�y�-l��}�tub��	x�K�����_�6f�lڴO������}MX��hHZ����}�E鈢ց���0�-��~�Y�׫m&e2���@��`��Ҩ���Ir3cʵW&%S7���E�	ܰf�hP~����=;w����.l��5�5m*��>�tqC �����׃W^{�#~�AH���S���)at�aRv���U�sAX��P�~Ըo���h���:�)@�l���u��k0w�����x�����	�`��Y�LZtE^nڴ	'N���=�����?0Ч�J����c����j�&2��F�Eʉn�o~o���~��5U��
��[Q���)���s��3o�D�)\u�5x��������	u�Mر�S��q������"0�{5C5:Ty\�����]�r9������ø������G(�¥W]��X�GO"�ʣ�u��%E�)��R)��/�~��_*��rH#P�n�+p�5W"�`$�B�H��<�VT�a,�0�1�y��~�Ga`�A&��wz8�1o�r�v��b¨`�պ�tc�;/�B�)�Ĵq����I�1a\��sh��#��&?	�^�c^�%�"���56������q��Y���FtI��q���Rd`F*�W��&���B41f���TQ/�ydT�@E�9f�R}Sk�?��_�����/~z��@���A*�G*�1{�h�����l�>�]��g�V��Q8,:I�3 #
������Uۤ��� ���ˠ��
��~� �ع[|�z�C�,����V'*�ꡳ�0/!�*IL8�l�R��p?��0t��(>���<�"iEAO�ÖJY�2q��15��ƀBFj�et�/���Y?���{7����D�������m��I�2cv�9�����T��K����r7ݸ7�������c�����zT�%
hnj�=�݇-�oŞ��R�on�֏�c0FN���T����#�1oH�
�Sn�L����)�X*"4:*'y�>�a����U�C�� �������Hr��/���	�)�$u��Rͥ�iP��6���̊\��+�u�#�д)ߧ6(����d`���Փ��a�h3˦�S�8q�L'L:��-�y���������{PYY!��];P��t�� ���]�x�l��.B�a�SQ��2��Q�Iϱ��P�#�bBϜ1��v��^�{�orO_��&�lزo�����XvI�p�5W�i�����WHg����`��ukn@mM�<K��,L��X
�r9�|�Zp�UWaђ�x�������8U�b��o�d]�É[o�sgϑM�3;w��^6-q�ׯ�ZN��Ǐb˖ͲH2���K.����dcOē8~�$�m߁d&+'H�i��qH ��f��ȷ��]6x�rV��-i�!���`֮:|��������q��ͬ=�K-Ľ�ݍ��������b0��҇T,��K�a�+E�����q�u����5Μ='ɭz�KE�k���2�PY8�w���#�2P����yP\�!��!͡�l�j�D�
8�����	��"�w���	�=NP#�	�#�!�&�g����I�g- �=b�$zz��5ӮE�M���Wm��x�;��{o���[6�g��k����
M��*��\�NcٲeXu͕x���D���?e�Q�����2¹��;����Hj�ʕ2b����v#�H��N��704��sx�pz*��?��`�W^��FF�
z�Z@� R&�H��L�}	��"H�G5"O�V�K\v�b���j�1�Yt��@��?Ni9�v�1�}
�v~�b�}\t�r��@�c�a���ᮬ�����,�t�$��h�@6�ֺJT��ECM5&L�IS��>FB MF��9u��� ���Y����#rPa<��W�|Ɉ��c(��h8_�D,��j�K&y s�,�+=0!'f�rp?�z�8�o��{�dg��*�K1�?�����~�k�F��_�+y8r��[�$��z�6$�@0�@?�iG�ᱺ>N���p��.�w�!���nD��
�X�h!n�~��;$��>�����OlGSKb1Z�
(���M��S<5pyk��58p�s���F�Fb"�Ja���t�*tY��$�s((�U▙���� ��iM�$C�%#X���95�F��M	��觹�
���
���q��	�67J�o ��
�g����S��˯a��O1<@GO��~�̚#�}"�5W]��o�	gO��g�]Hr���.�g�7�|��j{�������;8��;v�?��OUC�D%k��Yayh����7)�a��"�,vw��6�<�����M�J]C��.���Er�a�)'��򕎄c�{b�� �)T�s��f����/5.�g�\@Z�U�qW �y�VE��X^e)�"tI��J�L0h���h��45�ca�&�/fJ\�uhj�Ǟ�;��G[�E�JD0iRn��z�i$�a��jgfAV����{�ݍ��O�I�����kio�⭷��'�>��e�q�7�=��������臟[cm{��h�<��#V�`�{�I����S�z�Ea��2g���ӟ�,���W^���nO���w�ـW��7D��[ɤ��9�1��RW�b;Ȑ1|O�� @�.�R�����4��D��[JĘEy��P&9UJ������S��ی5!q��(�5�#���_�N����㿙�KfH6��/Ã���S&�G��{�a��F1���������s?vl�)�1�����QS_����/���D�cTO�J�ր҅�J1*�w��邯�"��Wl������gjT ��,	tʟM�zYft
�i�_3� jvz%�>��̿��*���`��� z%���z���O��7��
�L��RW��.^�I����04ЋI'��܅�[?DgO�0�g:�����ˋ-m�j���2^~�U?z�]z	��jQ]Y!�,�g᫨Ɲ�+���E��[�� 3N�����xy��8p���
Ԏ1�_�S��#|�����%	�Zy��pJ�
�����,ƕW�V4U��c$��P����.vi�H�y� ǁdD����5�aq�0y�T5�p������bl�q��d3�����n�%`L��b��ҋ/`��݋h<���.� ���o᫨���Ο�L⑨�w�m�1����.�CI"i�O����/GNoC�Ȩ�i6��8��e/Ȉ�9*9x}6�߷�;�a���%S}>�?���O>����>��|��౎�Ǣi}��S���5�\$��0�
PQv��$F������;�����hi����],�݇�����'b��?A4�¥K0i�d���94�5�����6��쨨iB$V�p8��P��1�Sy��v� �N�?ԋb*
c..�;|x�is>W4ڑ�S���R^��&�bO�r[�J��D޼�Jhn�C>���E�i1ᒋ���_}X���g��i1Ś��҆��q���������>TT����.��g͜+�Jpԏ��J\�b9-����0v��!L���
̹h��LڋϞ>��^~�D��/��gp��x����S1-�`Zi-c�#�y��L��p �S��5��� �A�L�%��q*,�}rY��ѫ�u� m.��3%ǘh-�������B�,��#��I�-�,B��@��.(j�$'�2�%Ӗm�e�a���X�ɞ0���02f�c��a��&;{r�������C~�+�����@_O�o��N��� t�,]43gL���d���i�e�r�L�HTĈE}]��~f̜�Sg��ͷ����B-_��R\~�J�54���ŗ֡�)��s{��o��[�9��� T;��d�����ÃW_}�l��/�m��*�?O�����D��^s=�j�"���?�����@�ٙ���+9&�zp^� �3�J�T������RfԘ���6�,d����6 �L���k+�mR��d�-�C��j͟!�g�X_�Y�.��&@���ve0U���0�R@
�N�ˣD7��#��j��$��8p�U����+�e=�ʈ�w��}x�7�%��{0�|B��cr�8w�l�*i��lUb�@ƅ`�|n�RX�Qn�U�1�g��� G\)*4Jm����1��.Z�����XIe=U���#�r%yJ��y%F��J�(?�����'�������hm������b���S��X�O����O���SgL�d��g����	1n�d4����;v�^��������\�J�n�X}{:;������%3��U�婐<�x��U׮��/��݇��s��k��N� Rc45z��2Pa�	?zɾ!P����cͪ�qݕWbh0�`8�Eo��xɅ�"@��m0����A������h?�̄��D�f��iV0#�������i���-�hJ('hln��X >KK-�@O7~���	X�nl������e&�E��E��=�tA�D΀�)�E�B��׾b:-�o�6�Y�Ӓ����Ç�PIS��p��@_HLo��������Pɤ�_9�1�h,��J6$2l��,P1�ĉ'�T�g���]�D��r�e�c1P_������f�ְ7� ��g���@4��;��R߈I'`����n�$Q[�&�[�HD4**}<)��J�@6@!@6}�<�&�v/�6Jz�8!����=���F%����I��VJ�,�+���	V����)/	�|���0w�L��2�����;.#Qlظo������'`����f�b���(Ɒ8/Ȫ��4���[>�h4,�CZ���8yZԃ���hq`�����39L�>S�E����o�ERf=���EGB����<~<z{zp��I���!����1��
��*�xr䜛����g��EQ�(|e�RF�Y䔬Ac�y����hQ��Uj� K��2T̿,�e˲V�P��Ǵ
�^´
�FH �4��g��80B�J0\�Y5j���tv�t� 4.��&Y�|����n7�|z���Ğ��垸h�l̜>YQ5��JϞ;�c���F
I��e�pz+��ǟ�����c��^t�E�q�M�4i^y�oxa݋R�'n���ַ�x�i[�{�P��ç��ܯ������c�Zl����)��w/.^,VZ�g�`������⥪b�OO�Y��IjY��4iw�E'��de��H �&�V�,te����S�b@�%E�XE�(Jf4�䯀�X�eġ��T*teӠh�������A���b	9�H�+d��m�R`ibΐ��(D��d�(vM��aS1���l�b0�\X8��{�� �!�R����,_v���X,���At0Z>��ϑ��$��:{!�(��aƘx�I�F�c��T�;��8&2�[�g�I�J[�`���[~-�����D����r�/`���j��#(j�4���&�u��E1*���;��.4�V�����m4�U���N�:+3�v��7�ҕ��k�!a�l�Μ����䙳��W���}���k�E+7`C�L�bC9��E�0�-��̵�Q�\ׯ��f<��U�;z�Dz���sܬt)*�Z\@������\g�4a�ǓQ���Xu�"�p��G"�8�E_���H�
�|�����wa����Q��*k�1a�,x*��&�]��Y���Jr�>������(�B���l�tut�Ӓ,���J�2�gu5����í"����$��.��ޞ~�� �c��4]��Ʌ�s.�KK$��	�?�>�f#lV����Q�s���v���S������
��鍕�������"G���H]6c{�t��뱬���EAgE<]����� �Q�<O/M����ƹ�`-��\]	���Ǌ�J'�f��Z��<Q����VBk�.����n;qLt��R�Ɠ�hnAg۱TUumHf8p�ñ,bY=��d��(��J��PJ���n�E���k��+[B՘�@��f����G��JZ������z��I���`7��<�و�˗aɂ����CUe��|��۰	�^~M����CCsv��+���K�e>24 �	�,�eW���M4�~�$�����a޹c7R�,**����ع� ��4�̚�������\%D�#�hΚ1E@��������T��VAo2�fJ��z��`P3t�ttw���C���k��\idN�YQ�2��T,�:i�Vn��y=>�)���	љ��Ӎvz'�XΆ*�S#��m��D�D�
7~a_��`6�*��E-imnll,�8� ?k����*	���r��;�u/�EpdP�[��k�rr�Ʌt@l��V��ʕW����w6nDWw/b	7�c���N�/�q'���;o��_g��~����C⢹��6<4 �ӎ��b�ֽ�������1�o۶m�*0������ߋN���K�-�{��_�yZ��iѦ����D.�t-�ڛ��I�!oUX��'RL�X:�d�'N:e	�Hz��W�$��N� ?GJ��2��<ԘA�:
�^�LL�^��XlfƸ���(��!%3Kk.\���\��\%Q�D��^���N�J�(�d¸a�y�oy?� j    IDATM���=�{$�(�RQ�C����Y����G���{T�ͽ�!�Ϙ�. +dT΃��23����ܘ����=��z��qM���2C�a�x^B��8�P S��$ޅwq9�"j��s�w��J-Mu����;�_Ƕ-[$w�����D<4":��� ����pi?#���ZEX}�ʫ����0���'X�~=^|�̛=���-d�R�J���$�H��I�6_���dRU7��[�����q*�i�k�1*
�i	�%�J�P���jn/	�b�+����"�,��P#I#"�\f�J�n��4�R
�D�XX�U�n1;�Kz��ࡓ��k��x,I��:���aL�ڎ�S\S��h ����H��IYΜ>�\:+)u���1?�����J�
��Ma��W�9��e�4��YI���<�Q�YwZ�Y
����k�A&��v���dc5H�Bzp�<��e��������/���o�?�;ǻ��E���S]�ߌ��Uw5�z+ `�_�l	z����;�ǩOw���a�lz�[�7�`��Ihk���� ��0~�t$�E�M� �h׌��^)��$������mZ�SQ�d�$:���8v:���)0�|ʩ�O���^w�E!:$)�e�-�Uv8+�avx��A	�*��R@%E����@	��q������I�5����u�b��c���M�
���'p��Й�hhl���F'�&��.^*��p ��!�#
��������cI'	B,|@YNUU]+���� �+HPo� �Q����j<�h�|mM�Lцʓ�ݡ�Z=7���y�/�P��)äH>`v��k�n9Y�f�Sm��7Ik�srr�
��ǨC���FV@�%kk��������3���l=�mi�S���#������t��IX����>ʺ�}�;/@j��E;��;�Mm��F1h�2����ɓ��X���?Ao�9ģ!�69VD��A	�ͭ�3g������@�`�[|���n�aɢE��;Dt���O���ϩHs�Mؑ�}�ۘ8���3��U� +�����=��R��~��4�>��C������0�쩨��#�<"�.,_���#a ��9��#N���[��*ԭ�*��# �n�jA|�s���S��������l?�r��tYʍq̢KfR��Q��H���tu夾�(�q��#�ω���6�<i�0LV��&�f����\�@uu<n�8�`���?0$���5�N�㫖猟7u2d�P,����u�����j.G�+��@�g�� 3	�,/�j���ȧ<�)��W�1��LY�R�*�;e�`�̠t�5��a��Fu=�E���!����)���,�ZJ9��6��?|ﾹ��&r����57`|k#�n;:;��$S�ף�Uu��TT���G,�K�^���O������)���/����ղE�1��M֮�
����q�o��XB�Ӷm��h�,ǭ�܋�x�9�=|�tN���&��J�H�m��
�R��X*�������.��W]���a"t���ֻِ���1�
0����f��z�v`���as��7�3�k���ݺlM�F�t���m�aȧ`�'�x��VzDW][#k�h8,�3�q>��4���Y!�r~ �{P2Ke��D�ϰ���)�0s�R��.�Y,JŃ俨�Y����i	l�=�@���]��E�k+#(�)$g�T��'���e������#�~�D�࣑���@���"��	t��?��7�7�`�:ęc�1��)�F\<ofLnǢ�31a|3�u��;�����@ ���X*�Y��	����#3�j_�V�R��m��݈����S���T�0]�
����9)���A��wb���X|.\x�A�N8����*��h�����L<�\&�R!-Uܜ�S�T[�5�>aOH��xd�Tx��a㰰�b�0�08��1����#�_�!����W���9|gO���g�Y��.Ϛ�ɣ"�3�Q�Ј�S��g`&�n�ݽ=�E��!�LDᲙ�ۤ{i����&�d�ex9�6�ʘ��*ֶ�؎�Y)����ٳ�.����p��1yh�Z�=!��䔳��� $M���Oi���u��������R�D��Z*�<�)ۧ�5g�J0U?[��,Փ�V���A��_���E�*XX�Fsv�(�Gb�ڴ>�P����H�l^F�gS�&0g�`�I�:
�8>�&��'�'���/
��4�g�E�f4c�����;0a|;Ξ9��gO��A'���"fϜ�S�OJ���|{���d����8x��0mt�P��o�l|o�ԲWVV�k�¬�s���,.F}������Q��(�Yh@E}����t��,��,��*3+�b��S��cIb�T3i��TΫ.�T�E塈(��Y�B^���A4��c��9¢p��<ׁ�����	��|�����e�!#��7��͖_�RR��� '۳]���M���4�O�|��1��1 QU����fp�'��|�Yj ���@���R�(�@E���1��_�a�m��rK��Zl�ҜPj�!ߏ���눮G�_�3h�Vϻ��둀2�	mM�o?�!�{����:	�#Ke5�1e�8�77
p�
��!��>�~�ߐ*�o}�I�Ba<������O�	�׿����L'���BX3���S�E�G�<^|�����/�Ok_ā#ǐe�59�6��γ1}�v͌D�ibZ�0�]���b�|��Y}=��G�8�C0eD��E�dGZ�z���Z�$$F��+�2e��U4$<P���Ή�c 
�0�+�0�����Gz�T��1��A�Nk[�0�tKRHƷ|����Eg��<�/��?��b�B	�T��E��[0�
4�O��?��@T��*���T�ag����<�lyv�L8��>�����M�\}ͥ���&߯���}�\ �Α��L���'���N���D�dE�b�PJ�J_0,}%�����E�y� z�D�U�yS�`�qX4o̟!��/����0f_�No-:�����|ǎ��U�����`2�E��euf��
c0���+����Z��<�ؤ�At��h�Y ��Z�}���'��8�l����	THu��	d��r�A��*����0�U��072/���몐#���K/4gΜW]2 ܬ�y�dٮ�ZE�Vل��"�p���/��6�*Aa"�-`���:��9�.��I�X� -v�����1e�8�Ty�u�,*�TWW��������R���yL��r��f�"��<\܀�<�g�}o�& ��"|3�(t�cF�6��k꘳�\	m�Z�.�&���\/G]K��E\:�LU�m9v\kD᭶�e��?�3
�0U�_��YEЋB��A�l�q�]v&;���sd�
7Y�z (e�HB]wjo2�J@`OQ�T�Z��n�|I����c.AV�N7�I�����I��h�?�<�̙���J�&�R�ڿ��$�i<��a1����2l.޲eN?.Y2�-�w܆�����tf<��:�޻OFa|o�<_#Y5����ʲC���Oى�Gk,�=�sQ#PQy�/��_�Ju2��5Γr--�M�d�H
�4��4wQbg�I̚5C�Z��Ϝ9#I��R�Df%�$�N,���R\	�lf8s'�%�nB��%�4��p���,�#G�PS%v��⒢���o�9���WL�H�3ԇzefeL��ٿ��9Pp�1��$���K�/�~�J4�X��bs��-��ŵ�À�I$=l��%׾ <��_J���0��T!���:���O�7��í[e�)e�����}n<n�=Ҽ��_P��d���5u�xi�k�=\�f\N���?#�QMס��|n)e.KT����3=�Ʊ`�Ÿ��{�v��8|�dm�)��q�޴�Gc�(��J-�Jfd�b�"�r�M�����aFK����ΆX���Q�7���Z>��4q3��шH(��4ɶ�ՔR�8J0�S8~`7N
}.�b*$�L"*�6�k�ݮ�Nl�v�%�=�L��7��p�SY�]{��2�,�M=��aʬ��4cJF��aq��}�g�S��JŨP���9]�YX��f=�O��y&�ۭ0�Bfxj��?�ڗ��tzs�o�������t�����.K�V2E3��"BL�Eo �B�4TXQ�y��N��TĴ�\4c
�/���s��������᳘8e�v��F�tF�H5s]����ͻH�Wc�&DRt��bp4�hXp�JX\Dh��X	�D=g�#8ЍTp��fr�V�?#`w�S� ��F��2G/e�|�@%��BW$�B+�yR��D<��4��Px���`�@�n`�V肸"8Sgo�*�㩔�vz�PVe���� 25��g��5!�6����3ɔ���ZI9�DD��͞蹎.I�4�-����@?Z�P_]�qmpۭ8��i��\�i�K�-��9S�p�db��/J��( �&�
��I�|f�Z���;"%�u"�q�<j��3n)���+��<����!��x�Hp�������Al�g�����kɿQz���ͨl�,*�	G��{񍰤��&�b�F\^�������x���m�\��V���Z �޲cB/%���)��h�#�&�R��I;$?�\./s�"�tG:����t��򢁩�x�RF�	i��X
3�Y/�A,FsK��A���~��a��B����hD4�:��z%#'��{�17],�T&����"L6�±���x��&Л��Sg���,)��Q���
(c�^�Po�?%;�Ĵd��B���ݎ�����m´=�� �I-����ļٳ�ر���ę�̿H/���[����@���M|N��E���@k[�l�̜�%R��,���a���"k�Ʊ�W)����T��s�Ţű�r;��9x����ˮ�rs���5����-��AJY�B�T[jV�2P�&M�	�t�8���H+���BZ1���6��Bt=Һ�X_�'��8ֿ��$��ZG�Ad�̑��lM�<��q*��EKhk/�!AF�6o��ȳ��?���d&��gB�ܸ�Z�c� �lɊ.Zz	��z;���::vF�C��2P.&���m�\MԪ�@I�%+k�KTcFW^�7�Y���8�IN�D0�!�sK{r����ft>*f�넪Q�:�#<��r�a�O��Y�F:��a2Qt�:����Lz��"��(=#��=O��!���h���MGW�0���>��tN��F�UM�5)\�:�F�fݍ�*%�����%�T���uQ�%�t)�ˈc*��`8��]pz,��������o>��ES����J�H]�Zyo�`��#�B���KV<UD4�F�2��1�Pr��"0p��?Eh�����&�k�î�M�A�Dc�xI�Kf��.�4�$ŒlʉX
��Z<��Cؾk'|z�X��Iؔ��(<�͘s�Hkt%�J&C"Blt ��A$�������Ab�]�jX\�[hg.��L>�|&�L9?���E
�HO��FA.�� V0�|rJ+�E�7oPnԌ�'=G��M�q�f��� �,T��,a^�.������3�+��j��l�#A��!{��(�����cp`@�.�5�܈������n�����Z9���oRJʪ6f3ȼEso�T���aEN�xzt���w��o��Iږ��l&/c�h$&��R�'c6%�!eu*��(D�����`>W�4:?�^��?Z��Jb�{�֢���b���l��~n�'����B\���X��볯��T�*��b�D�s�3���g�<�|G"!�Bs���� R	�TP����ʡtV�]S��9"����<�r��B;�h�̈�"p:�DR�U���EVD�q�_�t��M@,:��>�\p�vT��$�P^��\*��)���b�ZY���GYj	�T�57ޯbo�zmT4��4Ua[���(��r+4A-�5��·d�:�r|f�}ce�zN�M�?3�M������?�7��� D2��8jҀ$�+~��u�5��4��ŀ?(@�����bB��91ؐ ��?4(�̌Y0p��	��Zڞ�X�v1nj&�f���4�>�k��/��&l��"±?��ӈ'��L�G��M���V��~5���<�.^S�J�����P\@�.G�Z����jLdY/Cv��	w.�<��F�Lo��� �������
�O|�q�tua�3��gJ�U"F�ic��Sw'cCbW	�Ӊ��"�r�����$����xD��P3���T�s �Ԟ�!�N�WU��o�	m���wx
�#�Q�k%����Gǲ��}�ƭ�]P��Ku�Ɉ�/��7߆H4(����B$KVD3��YJ��/�i�ɦ(�rBRLf�BnjSd]��[� �����c1 ��Ź��8��0�8ZO�nщ�����{�]!���Cm`Um�0�oo܊p$��z��㦡�m7�єt�����+r]ˠ����z��4�Y�����c���	������������� ��,�FO��'�������VZeP �$� �� 6p����/���ca�`�s���@$W������3�s����f���[��e��]��t���9�	����޷r�ƾ��x�22��.5<o�]z�B���
��� _n`9W����X� �;��ʫ�]���#�;#Kz��E|�hOD�v���я���Ȕ
�ԫ�銣�Ϡ3Ѯܑ��e�[�׿�|��_ǑS��\�!Sn �e��}k�`�\6k��%��b�W2)�K9������E_.o@˥�	s6��'��艑E�]"*+ݓ�EE�1Q�N�����R ��g��!�n�NCH�y�Ysb�5�n#0�;jAyP�2�ɜ���W�y��/ù������$C�JE��ζ���[7����f��hH�/y�M�!N��
�3��.���Ak��-������w��=!-:h
e����sy]�Z�x�
��̖�cYCs�D�3srx����蠂��,��
�))$�_ݿ!��`6�Ӡ�<րؠ�z9�
����T�xl�ۃ��p�ג��s���_��yY��'h�&_=B��,��]�&���|~HXk�E$�RD$��._?y,(K�
���Y��9��x�5�����P*V������W���5�h����I�\u%F��2�# �����H�ϐRIR�!܅��1(S���OG��y�3!o�^�BU2`T=�q��Ϝ�9�I�w�����.R��SO�Zc >?��C˛�]%�*z�����,�&�����&�5"ؾu�17�7P��(��&��y!{]=B(�dLߣtzYE��J,�6?O�CFJf���{V�m�����&~+��"z��ra袊��>+��Va��l����Et�*L�|�Z�֞&�H���9����*%$��)�ř������ �Qe8�uE��q�m�b�e�3����l
L+T�i��l��+a�Z\Tj{{'�F��EXL� ���H�lxm���(�f��hokS�^6竇�D4�n�����8��xݪ"g��!��س��x~p\c#��j���cV�K��\y�x��oC2�E����L������BEh���Gʬi\�P���r��N��A�4��"pK✞�4"37f2��E8��t�y��᪄C:k��*5
��gRp���u��o6nۇ|��T�Tf�1}���*:�ÈX�PA?*�~�8u�����/���s�Via(���_����N*LOv6|o�]~�B���&Pm��+5��)ab.���"��Mâ���Z\���i��>�����:q�Ϻij�E4��u��[�&�T�m!����e��RNcV˿z�i�U,,Ps�����'�@��&��n:�:�K)�S*:\rګ�Y7���ON/j-�ԚE���V�Z��U���E�E�=k~�2�]�����d��pX�f!O��n�3V7i�y��	s	�����j�#8�0���Đ�Ve&�A7L��pRB�k"���&������U~O���Rx��OO �ܽ�z     IDAT��_r#������:�^A+��=�6�<ӵ�{�02sb"����8��o>����A��l'W�-�F�)(�D�\!+�!�����L���~���.Y��f�|����p3�Z�}��*�Ym͘����gA>��!��qL��5�e���ݞH(n����ZGO��h�L�%����gb�*(-Vv��3�,���Fб����It�v�}�D����GQ�������fC�.�|����[�%G�&��s���B�`�a�s>�+&����w��������g��X,�`<X9~�/(h�2�2��K�x�xk�%��aEE�=͈C[H�Lۼ͌�X��9h��e�o�s۔��k�]������_r3�F��?��xml
Xl�Nc�P�u���юLvIH-�h��M�4p��CZ��ݧb��j���
�&'�t�2=��S$�*U�E'���X�0��sV�|�F����i��Tֈ��oI�-�8�\f�Y��J�`��
O���b��wh��1|#0�G��N{/d�b"t*��%�!���.�RDD,"��e�HL��Kr��7wlۊ�w��"�ըVb
;�n��A#����e������f\q=n���
��f�BیpF���9Ј�����.T�87>��Բ!̯����K �y.&��1���E+N�id˔c��2���Waj6�Z+�����(#��'��lz��݂�y��^")�1`�B
Z^(���,���p�z�4QX����q,�O�ZX�2�8�e��Z�%r���y�(j�Fb��F:�ub��ź11�D�T���ɩ���V5��h�-D� �,�(���8{�Ύ�C����jV�k�|��?x���臅��x�����Pq��Qi���װ�)*�2�)H��l1��mI�e,Ώa��$'ǁr��z�|p#NN�����&�Bسk;�;f����挳�8v��~?�ŊTG���[�g�5(�]�W$Hc,>�l:�lz�j	�FY��P�67��$�Q�1��p8���U�T+��4�3D�t���Ɨ�_ArH!���Z��C����6�]ٮ�������y����qxᓳ\u�V��#5����qu,��Y���=#7��7b��*$�����d[��7� ؇R�*x>���BE/�݊�c�<��F5�{8��������c�F�?awDE��|��*�L�a���]����ֳ�/K���۱.[�zub4�"rS����s��ت^F\[�L��{�e���$�I9<nڴ�pL�%�D�xqQ�@D��.;
V|���(�V�F/��B� 0@Ͽ�k���%�SgQ���3y���s��"~��#�cL�8w�����$H>\N-`fzܘ�|"ў8}J���-�Q�;U�����(�zV\7���K�F�Xp-���؎�&;N�+��m���`�t�z͚��b�F����֯�����m8*����w,'cYǓ�C��r=�󕷣�=�/|��0z���|J��7���A�z#�؋�<N�;���ˮ�\�s�ݨvb4��ҧԛ(	�s��8q���)p
���l���T(UPUȩI�?�37H�w�8���l���*����X5˿F����m>�1"4kD�`�tl���uT���I�y�<d,��#���TF֟� �ǋ
��M=�R!o��ؓ>�#��[QM]��٘S��b���V��v�~	h�O{�[.��k�g�C��76 \v|�,�X�4k55��n�q����V8,�5�0��(ך*��9��*ޘU�|FvA�B��� �B@-��
6x��^t͵��Uwadt��禳�ɢ���r��6M�J�hq�y�>y����b�2����H�#�>UC�I�](/���0�����4
�e�c�,5�B�L�!� ����c�~�����(@�r6���Lp3_��B% �5$x�TB:��\�;#÷}���y]�YX�������?��'ӲPi�|o��Y~�B�����L�B%���,p9_D�Y?-�~看�I1����S��Gna�ZF���Eh�	��MN�%��?���K/���$��<֮ۈ����w�~�裨���9�]ု��_y#��>���Ĺ�yHs������*��`
��\��>�k}#y�Y-�Vf�OF�E��M��|��*�%"r�e��Ba_�I^�<4�a�(�إ-3j�EW�B&���&�~!Q�3]	BY����^���.z+���Ī,/�qsN|Ӌ���];�����YEG{�3x�o���A˧�i潙z�X��'5gN�)ΠU\Q��\�`�b=���/��S�"�uuv��gF�< ��kq�����a��yV��s���V�Rq�Y��Yq�����P�Cc#���lݲ'���*o@��]w݅�T
���7��p\�K�L���.}~+��!�v,�"��8�ey���r�W+��h/�g�H�?��O�t�ر��Y��l��
� E��YK�� ��F$Do���P.dU����*آ����+
U,r\�l$7����LDSC��
W�O8��ǌ�b�$.Q�R�s����O�@M�=e.RsގA����3�a��״¡0D�]rVL7o>g^�ձXBK�o�'/����������)I�%r�}D��ܦ,y>T�9�pw�%�&�y���8�FǕ��{�N%N���2O�����9>���9K�Rbp�V��g.��+ln������W��ϧ:�(��a���tdS���*���[�c
�=U'E*#=o� cH�ܵ��X���9��MW�R��{ۨ�������X�(�u�3*�XH���/�?#^fD7�V��#�V&ycu{b����!��dٯ���u��{!���s\�|�Dp�V$*(M'�% D�(������C��mH�N�f��c�-�8ǎ6�'�E�Zc�H4�cH"�lrn��%��N����r�&�Pn��t�T���j�:?��`��P@zp-�Ϯ*��b3jL2�d����!/-�ɑ	��E��M��$��R"�D�hyOt"iC��q�je�8=A����CE�Q��D��	���B%����4kJ�w�X���tr%^��<� O����/�����m���)TZu����3�Y�6U�Ԛ^,�kr����W�GD��0
\P>W��r�y��:���8��Y�]U4�YU�oH�"P�FU&B�kU��������gqvbZ ;<p�;0�n'��\,-�O��v%�aڒ\�F$��͸�4��L��Iʑk��Ɉ�B�A�
�"�()f�`�==�{�*FX�pS�a��ۣN�04M����9����8D&8�	j�>��Aś�K�G-�,�l��6AK�f$I�
�
�ёs��K���v��زn-�G���[m� n��VD�͉�>SX�cB�+s���n��Gn�VI=�%�0FmA�N��H����?Ʒ��=�vƢq%��p��8�^�"͆�S)���Cr�u����OT����mm1|�#�?HGg��zJs<Xy@s��C���Pyի^�C�����Eߟ]�����ƙ4G0�{Wu%�:����T�UUhѸ�n�j-�{U��	��F]�2�p]�|K���F F���r!��f��<�t���\��h�N�OO�^."�qcnnJ���5C��ې�Դ��RH.fQwxQiP�2<+�SN��d�Z��x}}��,O�:���9��	�q���:�GT[pli!6�D�����(��/�* G[����a�L���r����^��;0?7��~�!\&Sˁ��%u��v����{�Od�E�&�O�`gF�(����.V6�-e��ʫ���-�ݟ���OÄ�\fI�*U"��p���[�*�ޱc�f�*UV '�{b�+�²ާ]����t��˘�BTt�X!��W���GMT X)�^mgY����
v�V�i7v!�����,�ju&0�X$Z].�%6�4�������P@��M�q�6ʴF�L��K��iL�(��rC��N�Z�6�ɘ�<��� �N�|_�|N�?#�\ҹ��P��lXl�'W�pH�B� ��:�p�%ߌ$W��`�O���m{Q�9�~�>8�=8;��B�o�M~%�M!&d�2ңJ<9dN����w�*��֒�T65%�󭳐�]J/�N��@����A8���0�ޅ9��^5T,F���{�����4�h��Qe��4���(��(sH����]F�<�P���bjK�#���o��%������x��ɼk�?)T�ȮΗD��MF�T#���w�Y����Y̌���G�����B�BS'2���������R��P��4K�z�`P�3��o��M{��P�:K�C�9�bo9�ZLbqq�؆QN�(K�i�y�D�xA�B��Zyɐi�Ơ��XH�0�l*��Pr4V�o+Hxd1B'Kn@��KY]�h�â��+�H(���vbq)�0;�<xu�ԭ��f�R�X*+_%6�/5��&���:s����f��=�عk+���Fz�s�P$J�W�b�"�c�~K,{���V�
�$M�`D6�7��o�W���γ��m&J@�p��9��5�R{	'�Rʮ���(Ft��"Ȣ���B���q�Tŉӧ���L��js�d��/~�q�x��ʽ�&��"J� F)L�&��-�ǆ�U𻚈����R�a
s�c��~����2=�<�:��*���%��Z���5���e�G2�(��oh�O��x0����Fqys�*�R�8q���ޅ��~��E$3E�᱐�_B�/���Ⱥ��[�q�\�荿�����-۱y�6y�<��Ad��I��P!a����Q�u�	b��B��S�h���Ud��L�O�!L�Bߋ�M]��p���`߮����F~y	�lZY1�ݝ8u�9�!l۶]�#� �U}��H �t
'O���j�����j��
�dҋB\I�}���8w�5�u�ks�Bi:���0�5�L1�Q�,(,�Z[}r�͌r���nh�<mTC͈�kv�懅(�K�Ԍ:2��0Hk&�I~�K6P$�Z�uOٗ�u�ۯ����y���|w�N��D���
�9Ż��Kf�D�*���1X�d���*�5"@�l^�-��sQ���	��ƌ��#^"��,����$ʑ�I)�b)�U�ҵMY|p��l�Xն~0��N�}^�K|-t]5�??��u�*�7H�)��^L&Q:3z�E;�����гz+F������	��T*��:5�R�ǙN�X��b�"����JC`�<��ߌG; ��2M��B!�����,�R�fˡ�])W�Ng���z�h����zѹN�>%�S��Q��}�	*�NQiօ�d�)�ӳȕ�h����CB����ց����Mo������f���7��e�0�it������#�� *�<�<�g�JE�Ĕ,�`�|f	���'� ��,9%!C2L'UQ�@��w�,":V�-��!4\���t��w�0�7"�և|�G�UE���,�D�=����Y�AB�+N��d�fb�cĤ��/��	��~�Xq�gHL�`P�t�8m��X��
���r��;Z��A�S��.�2	ۺk������Z��<�̙�kx���)W���Eiք���f�	1<�Z3�K��Aw""�N��4p�uWbph �X�bA�"u��eG~Nk�lp���,���,��)et��mbloxÛp��i�~Z$��0�[0#2<�̌ڋ��������%N�ɠ�-4��n��6�e��1|1�+JaD�ƌ'�x�\�n�r�-xꩧ035k�RY�z:��.�T��"!�⒝��g(	��t���΍� [,iiK�Pd G!��z��HM�*���S8����Q���P�W����8z�^'�������|>/���/������S8z�0��סo�^?�E�N�ctzK�*�-7\ްF�]�����bN�h�P�u�Z-�-[���ަ(��}����S�#�+�#A��N�ȵ��sm�"� �̜����Bs8+H��Rs:��,�M���@i2���"�n:����׽�Sx�೘�CW"�B�E߶m�0?7�C��T(㦛n7�J�[h�������y�ulX�A�|f/6���?��8��3���H�|��Y)W����Cp�(�.#�!�2c����ߊm��6M���&�Xo�/2��+�q��x���/�h�h
]�J����e�����G<r�*�V�g�Q��`�P���5ezhbG*R*����+�k�gH.�o��!gDb�I27�D�X�~��s(֘���.�5+r�6v�p�x�����
ךy�$˛�ʆF�lF�}X\�����K��R!�wY Qi�k!2��q�<}�yi��X%��Q^UD�3���#~-�*u�[^l�u9�6�C:�D!��Q�������l�2e9�ʎ��R!��è���O�J��'�K����ʈ�0 �\	:�5n#d�>TN�p�0�粱SɊ� GoY.�j�z�"N�Ϫ�N5��Q��2�X^^��9W*��� Xp�����}o�gƗ����������d���wb.��t�����%��pn>���ʥ�>H-X]3\x�0�xP�Ѭ���$�0;���Q�rꌙ��6f�l�����<"(A�toމ�ፈ����	֪�����,i�ȗnmՐL� �]�!h+���b��������:���i�Q*,�RX�
�����*Hܢ�[gG�:.^`�xB�R.�E��3C_ʪP���eM�%�r�,���f8�X#NNraβX��IR��N^�BՔH�օ͟�5��vQ^v_�
:�����8������n��t�qL@��_�^�=@,��9|�����~�0�u��[M�~����s|��_�X+�"�֡�937��edt5�)x0���`Q�.7JY^y����H4L������ad�uO�+{|!��:��\���Ϛ]7(�J���������13I�x��KHvա^* p#�Y@W'��[��[6�ת"�b�Y��ٔ�d|z
�̒f��^�Db/��~�	�?zJ�G|�uGk�oA|U7��U�e9q�?�$�L~=p�e���穯�S#ŉ���l��>2rN�ŗ�G����삊z�����ˋ���B�����"bF������u^���_��\�,��?�����q��\'�~�v���\rUH �o�]l�_4�2�z��������H`و��3u��L�n�m��k���~|��q��)��u�Cr=M��T��l�{r6�����I_~���"X�j���H�2��X��!k����B<Y��*�P��&���|J�� ј�*A��9m�^���:�f�Z�!{Ϩ�_1y;/a�ЉVE3󕬋T�Y[�<焿g�1���?�n��l�tVD#�\�zq����>��Z��\�A_P�T���q�:��(�c͍7������T�I��J^��������h�HD�%Itfz!��{w�Q%{v(N���P��qK�X�\>!+T�p������$��:�:�BWw�ۋp$��M:_�A�1�]2*u�."�|N$�3��_�艣�e�k���[6K�ε�MdD����>_;�B��@����U�_��X���4��l�hB�R���Y���#)�B���שD�b�4�g�����
m�R�c�&�����anH1i�3�&�RAE?WfZ%�F����<���q�s�	 ����F8v�(d��*S����92.!_* �YF�\D�ܭ�>W>G)9���������;Q���n����B��H�P�&{vn�$J�h�e��tː��0����䜭�˅FlI,&�4{.��Ũp$T5�v��P�Pݽ��ބP�C)�5:�Q*�4A��j�lf��
��d3iY�+��i�Tv�".�b�ƅU��р�UE1�B�����&t��T��p��i�����.���d�"�1>�n��ޮ^����w:+Y��\3��l1�����GD��)�R9!�)7��.�6�����ѡK�R.:`�p�2�* ����WߡQ��̘$v�q���;�f�j���4���r�OU�r����e�v����@d�j��ⳟ����h�J��f��F�������$��X�i��UE    IDAT�����v�$��u����1�,7�!�f�g�N��δ#��hKt( -�TUy9y.Q�_=��H��OY�(X�&U:<fp��ah5֯^���� �w#�Q)���rH��\)�Ny&M���?F8C��A�'���$��@�I�*�:��܊�P?2T��8z�,~�q��� z�u��%4L���L��h�x��&�u�^|���Ec�O�05�(ʹ��#_�!�*d���TS�z�ˍu�ø��+�z��ݧ<�o���8|z>+�f�p������Ȉ�$WT+�/�^�f���l��W���*\�=����.ݷ�\u ?�g"��N���K.O����]#gG�a2$t���2�W�P�`d��2XcZ�D]~��_�С�jHȿи�EI�(�k(����1��o%?��9�~֛�Fe�>��_6��H��w,u�N�t_a�	��b�B��`:���eT�2��K^r���m����+����9=vZ3��D�K���y��ɅE|�_EWo����i�)���ł�Պd���bQK��p,
�߃r��L����կq��9���w���W���M+���I8F���/�tv$:E�O��ğ�u$T87=N;q���q�޳;v�T�@%���������2M�>���2~�$�����ϟ�g���t�.�L�$E �FI�k���y{WN�2%L/06��\Չp[]=R���Y����e�XA)�E�G������|��|�`T
>��x���P�Z�\��V
�
!���]Ad��D�Z����
�~UŒ��W�P�-6��AD���Y~DߨS\LS�R�su��V�b���Y��ULv����m��;Q����u��7��,�Q:���ۑ-9�+ք���/"�g���M-v��Y�@�k�#�aQª�P��e�%W*T
+�c$U�7]C�]��k�13r�a�|�E1P�!��R>$��N-�ci��h�Ym�'*Ɵ�
��/Hn���$\WD�@�|y�Pa!�7g�4üL;;�`8�Ⱕ��1��l7� $Br�⤔�T-��ץ���ng��a:(��c��P8]���l��H�!N�uS�3Bx�` =�m�x��/C�\���5��������6t�v��ł�B�1��:�.�fѓ�-���lnYőפ̺���ѻ���hIX�:�x��>{�ݽ��'026�N=��%$%��F�J�X�����z���;ё�*T�iԴ��F�az����-�A�<�����h�lG,ކ��\qi�a{��z�����#
��IU��~��Go"�=芆��Y.�C��p3���Y�l���ۇOˣ�}����um݄����8��ۅc������Ihf2kOw'<`x��N��(*����m_z�$�{1�)���F�搫4��˼���Kp����s�����h����kt�:<>�b	�Z-<���8tj����FYQ��������O~e�ð-�eQs���no���_[�e�� �}Lh�t?�E��oB"�#�T�W*�H0ް~�oϾ}��2��}a>��Ǐ�ꫮĎm�U�p?����x6O����>t"',�Y����ù�SRq�a�ى��ヅ
e�^nI��6�N�#鼁��3d.� �R�XÌ/����b�fm5����^d!c}���㩎;�[6o��'D�&*�3$��1}8*�F���8F��- &��Bj9��U����;�E��Ϝ9��L]�:��Cil�^R���Xq��H�;9$�z����˯mrj<�#,$礤#Y��A><�X�,��+#6b�zU��D/}�-X=<����O>�$����%J��'�i7`�P`0�l>�"�-��[�m�8�{��~��VY"�x$*$�V�A�A�Q�7�ŕR�O�������K��ӏJ��t�'���w�9rj@Y8ɹi�F>#��������Q<��l3D�~_�M�<��!���~�����mJ�PYCD�)�����F[�A��"r����hD�}Dl�K9�MN���W�9�XPp��"L�-�,T��ݡ��;���ߙB%Sw�ydf��yt��]ȕ�����Kca1�Y�{U��9��%�V^�T��9lq�8��a΅	A�¦l�t�$m1�Y��u@�&7��/��FLToв�,jk�.ϋr��K"�rC1/DP#=ؑ( �*V��c���g(!�'saQQ����a�c�;�W
c�f�i�t�>�����.�� B:_�M���b~!i�A|. �����Y�Ģmg�U���TW5Az�-��AD�.��{���<���W��������k�a��Q��m�)̸��b�&���*"�Zϓ%?7���,��:x�:�]
�#�cfv^��,>'���G��h�ȋ�ai�O�</�k����/A[,/gC3���y_��7q��1����B4���]=�z�����d�dr�B}6쾼���n'ڣA����OW<G��"}`*��hh]�.̥RX���� ��E�çB��s��*Ӛک�O���X�}�?t:p��Y��Jb�D�oBoW���7�[�J.���q��K8v�0��K�w�_y5b��Z����Q�L͡Tw�J mW��7�n)�Fr�R�:b���������#�r&����,NM�"/{x��YI�2��F>vF�u��hߐ�VR�W�����fx��Ì����H�u�b%�╷�.�ړ�=���P���>u�T�9��'�����a1�R���/�����σ��$���Y��a����}��Q<��O����!����\J�XL�@J��KY4���D��G�Y�.0h��35B��4�[�Y��v�U�,�hpM�����X[���9sV����|'�{�y<�����a�(|"�&�a��"!�{qZD�5g3OeF,"\z� ���?Ĺ�1|�>��Ƒ./F��䧐�O����HDo�>,F]f���Y�����غ}����B�@�Ԑ8��;>Qzr�p�Q(G|�e�m'��Yb�T�u7܈��|%�������d�ae�U�ӡ�c�D���.�)�k��R:��?h����� F����OZ���GEl��:J�g�'/,��\~e�,f˘Mf���j�����C��S�I��sָ�+ă\��|Tؘ�:�xTl�Q�f�r�mko�j�� �w��#�?&gd~�<�E<o������te����<���{pՁ&H^Rn�C<��q�����3�����g�}}==x��n�К�I?�_��פ&��Pi:]���PA�Y^X��������y�|w����l�K%gg0ڍ|م|����%,��䓡�B��t��b��'�,8JΫ"�ZNxu�ӌ~_J�W��X�Р�e��2;�̕�19-��Xhr,-V�c!5/���/��7�D��f:
�������E��a W�b4��d�G�_G"���C��M���)���`���"��]n���b�P�)�D]ȫ�;OΒ�'�M`4��J�^e&��$b�y��8��VЕ����/}ѵz�8r�9�0`׎-���t�q���ӜR�7�.,V~[�l����g�ˏ_�����_��_bddL@"K��ց����|D��&�V�_469a�
��5YM��~ݫ_%�/Ѽ�B���m��� �=�8f�R ��.{jv˙���-�9w&E)y��m��9u�T<�Y(�S�SU���E�y��M`U"�f�ru��Y>�:u���),d������Etz�;�tn��|�J^�uGC�6aͮm�y�*V�=y���OQ(�����[��Byú5(f�0C��lG��RjA2��W]+9��bgƦprl�\E�4F䌌�m�a��R��3/��(:;���&���Յl��љ$N�O#Cx�5��l�_���$6s�Z�&+`2�(C�����]\&r���g(���πϋ;n}9������b*���}ظn��f���s���!X���}X�zP!�lr�Oy~���'%O���Y��7T7rm�94�?����F�؇M��@X�B6_F�P�@>2�으��?+��]�[�&�P�3�@1��v�y��m�o0�}X,�l��=؍ m�uȱ��u��׾�5����Q�2d\��uÃX�ץs�� ��|4Nn6���A��������O����G?�O��N�!	��&�bQ1б^U
{�
��:N���'g�=CO������{�~|�o�^|��USU��cㆵ�!�p�H`��d�Y�`9�sc;lڶ�~����w��c�O�P��jh�X���7���KNʼXP�H�3+����?S�������l�}�3F�W��zZ��x,�M�����$_�,c+��=��'Ρ�@@�x�넪��ك��a�@r9�]�Ά���v�R6�V���&'�193��v�\�ދ/���߉���L���Ry�91<8����&�NO���֘��i��[�Y�D�X�0R�cN���r�O��������u�f������ˋ~�����Te>�C<�`4��Ӌ}n��E�YE�YIwF>��7��߉�dʓ�Ǜ&��J�]�P�$s����Ԣ��<�ϝ>��F�A�V�"�ن\�rp��$=����8/[!�Q�O�y���\A.�4�҆��J��t�aK�|��A;�|I�T;��v	�/\qTl����z9�j9+�7:24��ג�Zy<~�O�m\�s�z�+��im��Q� ���a�~�@�5a��Dx������g�AsȔ�r������|�8�*��XdL4X�߇Mk�`�� z;bHNN5�}*j�z�=��nG�ȃ��2��-��^2v^���%ȊǆL����H&�	����v���?��_wvt�N!E���D�J��z�V#W(abr^^
$��F��0<�[_v�z��*R�)r}fp��Y;v�<PH{~~�W��v>z'O��,՘�(�X�3I�y�kI,#z���N͚R�;"A�K���c����Qͦ5���:�n���dz�a^7m��� D�䯞���܁���5[7ap�V�n<n<q���#*�xp�7chu�8FÃ�P��05~F|�ӧ�azb]}�p�eW��K�36�±�#�[F�Ԃ�@�|��4.t�C���B<�$���w� ��6���Yd�&��A�.J�<����<����3�|�էAYM� &�7��,T�D�ݯy�x5GD)�A{[L��rZ�h����N-*M�* ��m�.-:�U](��a�3�m6�{\��n�y���Q�/��_��\�����G�L+�[H��X�T�����<�e4f�2��ؿg,󩄴�E�iF�*�k��yދ�����H�]���h5�c�6!�_��p��q!L�N�c��jǺ��r��T�(3B��R,�h��g�Z"Y|�X;��G��gF�/}Eɟ<��{��p���ω�Z��Q���YŚ����8z\���o,����X5����Obbz���4j��H�7ц�5�Eh���TDeLz2���.�����U��M��>>��O�Бc�S����������}B����֞x�1֣c8}vѶ���9N�&q����32�������^�t�1��-�J!�BH�m�.�u��� ���c�~�r���k�����-�f��N�v%���G�L�|FJ"�H�u��7��#=�����SX�qn~٭��w�G&WPlE��7a����ډ���8s����';����鵯����F�'ikp�c(�j���{q��_�-[6���S��W���.�w�v#f�|��_�g�7)�Q�H�
�K���|:�;˩5������������ꇡ���S���%t1=9S�J�27�����?�4��D�%l�g�c!���̔�Ͱ�:eH��޸�X��182�i��/��!i6��.���x�2���GhC>[P5�L��2♈`����Z4j2^�*�jn':}r�RZI-�b!���ݡ�3ú��4�:�$���.f���gB8V��p6Hu��H8�����S6>������ǂ׽̸aBi���ϣB�I�C��^ݏ�گ(�h8D���/�/��z��0H]�6��Z�o��4�F]C7�0E+o.<���x���m"�$�Ai�@9�E��n?����fd�R���,�]v!ʚ�l\�W]y�:�096�ɩ1���!�~&��t�Sz�vG�N��|���;4�?q�����B�I�B�����w���`�+�����]�3d����!_����\UMԋ�G�ц��$N<�,|�^u�����ݴŀ%��>r���(�HDt��W_��CCz���nS"���Y�^�'�q��Y�uva�9}Hf��O���1�,PsQgv�,�:/wF�2�����EZ�Ef�^��Lj˕:
J5��=�e������V����Ϡy��T�ɳD��X���Ϻ�%�(�9q�+nW��r*������"z#m'�$�c���oߺa����L�X�����}\t�E����!	pm��p!�C�[��ǧ?�i<����<e|४�6�nu�\���Q�J��X&n��8_���b�P�'b+�B:ۑ�v+�9=6�b7	D�.�� ߄g��]�������8}��\&�vv`��a�t�c9��B.kPk��Ke�]�v����O���s4c����?q_���U�P����c�t�'�B��`���V�A��3�'�-�w�4J��]�K�w��_}�C��r��`MO7���d?@��)��08�Y���qI���=u�ylݶ����ۿ�0Ξ7*�fk�{�q��FJ5:�;�BvX�qT���ĕ�YQ(�095'�=�}���������X���`_z;��lհ8?�X̯(z�X�#ngW��{��s/���,^r����Ǉ?�1,�3:�Y��BwB��Z)�R1�b�#"�<�8rd�A�������k�ß<��RV�tޟ�7myxÆu���bz��u���9yÍ/�+_�
D�����Z�ܼ�z�#c���k�׼����c���K�iK?}�|���t2m,AH�.� ��5���PA�QZ�|���|�?�NpT���wr��N-�� Srt9�	�J@�
�%���Z+��s�>���1����aMo�t�׀��\�
'���i���&�S���I��m�i�ۀ��Z���%�# w�XA��~lذEHCv� nQI�j$�Um��L�gt��_�R�4�Ry4�Ek�԰P��ʃ���Ñ�V�̏�ɼ�iP!��pX�υ�$�K�*\V��ȇ#�L��0mKlZ�����L��/XvyI�%j��`�B�$���\�&Qx$@�~*~��w��V���EҨʱ�Q�/��b�������D��ATȺ�/%���Sg銹"��^<��c�@YL���[5��ҙd
�x�V���e��+��K�H ��Vﳅ���08�gr^R�"�������B:E��fMRJ����/���9{
�N�4]�œ��\�zIc���6��ö�UX���C�O�rAd��d
<8hE���G0B�~?�� b�0���O<�#�����;�9<��ǁ�ׇ����9j$�ܸ���B��. �I��x؇�Ԃ.�p<�[v�Xf���Y�ى9d�-d�$�1���h��l�R�ú��=gry��	��p� �AT�@BlC����g��ȶ��PY�[��r��}咶UC�Q#����C�{����ضi��e8��X��.������ڍU�}"R�������
".v��=L���,f��ӟϦŝx����3���%s��8K.������B�ε�<��?V`�]��X,/)�;ÂE�xV��q?5�X�|��-c^�1#Q�lk[U��٠`������k^�*|��_ñ��Ȯ��={d\�0=5�TrN��l�r�,zzz�P
y���!������߃c'����yu��b˦�����䱣J4���QG�QC��	L������h˥*6l߉5�����Hg�%}ե���#]V+ey,q�ͦK�5���A�}�=�xG'���x������u<��a9\�۵��m��H�(-,/-ȷ��c� D�-��    IDAT2jܰi撋8|�^���0�L�߿��۷mQ��yP-�Ѭ$]�S����S|�'.e�h��k�sbd�6mê�!|���c3B��>p�:bȧ�Q)f��A��ղ�%�sf�'лj��؍�C���eW^�/}�8unT�󍛶�Mo~�FP,�=^s_r=����?��)V����E���k�R#��_?��}�s*���}��C�yV��l����g���G��B�G;�jZ@�[�A�N�<�'�B���ڮ�G��η|⚡6&���?�[}T�����t��
�:*TH⛞Mi�X�d$5~�׿Fzj�'P-���a>e=N*�#Z�29��Z���2J�AX<��#@�$�fM	_�V�l`~H����Wb떝r��f�?��"$�?�P��W��5����Q��r^��;�0��0��l X� G��n�J)P���EF�z�lC�au�DNX�lX�^R�Tr�#�իW��ra||�Z]�K"��R���רK���`91���s#�TB0���QC�G�~Mћo�NFfm� ��16rZ����Z�۳�XH_�f�Ae�d�f�ed�5�~q����Fl2֛��w��m�w�}B�x֪���004�Yr!-����v"�+��s�#��$�H���_߃ߏd8��xp%���jO�FK�A�h�eg;E`6��E+oDfJr�d���M7ވ��	|�Y���g�z��B��.�F���h�����c�P?�b�6�piks���O �ɫ+c�y$��֙��� �`�FlGO���;.����D;�r�4�x��Q���g�l�#�j��~9'y��qaan
�PP�o�c����o`-���r�Ne1:�D��E��9�.~~42	�.I��<x�{�Lw�YC�� nJ4�"a�RP�����rW����(׽�3Mk���8����BK�Ff�H�`{��ԛ�����[�q�0Μ8���NĢA,-.`~~V�7�<�ktvt`x͐�v"�h�=�Ẵ����L�'����r�ɥڊN�SS���'>���15VTĄ�1!��J��9�h�V�<����p,�٤�KM3�f���r�PY���c2�	�z��[#"�q[�!���.������+=��=;���_��|�x���Y_��شn-&'F	�01v3ӓ�����E�z�8|�<��s�w�%H.e���Kq��1<��#*n/�w	.��b�����9#�-� wK�D�]q���}�lشU��m��ؼ���aljZ*���~P+�̱�ۅ��Y�7pd�5D����������.L����n�W��-<���Fcس}��:�D�i�����H�T����9�D�@ 9@ƿQ���8x�8���Fq���#��ݲy#�_||.:�fED���D��H7��ՃK���aÖ��4"�@U�?�	��&e7pË_�j1�xȇ�xHy=ʝk6Q�c�G�������GN�ťW^���3ȕ*"t'�:p��W��*Y}��-j���*��=z����M[[���ظn���������=��c�^�6w�}��_é�I8�lj@�tgv��ֺ�t�ܫPȍ�8*�š��#x�[>�om����J��7,,Wޝ)���0r%2�F�gĤ.f3�؟>~�3S*�`�;]�V�l����y���8��k`��q&5~T!��Y�f̣xT��턗�oz֬ö��T]�se���'��OuF�ۅ��U�a ,�	��ڨʕ����QC(�C.��|���� 	�աh�ʊU;�^�DHZ����8�/f�t��)�K�%y,���eM����(JDr�N(�(�f+��"�ٹ�<�%I[��^�=�.�d�W�F[, �Ӊ��y�+�'�4��]��?��B�j5K]`]:V@�����h[OnK&�tɠ������B<�8�u1��p2��]�^��ύ�aW��p,�^t"f��e
�-�VAz�>4�_�L���F�#"P�ȱ�*^�I.��\ySx�'4V���U����>kJ�#~7�b���1�<-x�uT�y�+%=~J!��8H��Q��H��S3�<=&[o�5��ֽ���G��4�����g��s�����ݶi��L�}=�C�OO"a)�/�R�ށ5X*U1��(�s>�E�@��d�Mb�eP���sS]*iL�DgƼs#�X�r�A�C����j��j��tV�K�K�"�ɰ��\ol.���N���������lV�g����	�tF\�g7voߊtr^��CkV�_��cظq���ٙitutb��uFn\�k�A�	�����F�_�T5�Y�U�n^�\����r$:��f�O>�A��������ղH%��
^Z�;�,�In'�"7_r�X����\�\�r���"�����A����B8y�أW�u�TRmS)`��x��݅��g���������]�U}=��_�G?���
��~�T�#�7d�?���c��Y��_aӶ�X`�r�e8|�8����u��۵�]}�ss:[�ҋ8|�9S�֫p��R��t?�>p%���o����p�D;�mߍ?������TZ���v���!_����G���^�ܱ@&z��⹃�P�Tпf-F'�q�-��7��=���_Hizˍ7�3�E[ԯ�qr�J�e�j��!n�]�^��\�o0���9��o�	�l���O�y\z�>�A�����E>���Ԙ8R��M���ضu;R����K±vɟ��?���	�����44(���$��0:=�B�vl�sbh�f	G��˸憗��?�	���
�����<p9��8u�P��TSv��^�U�T�Ϋڻw��%��/�/~E��k��/��vD�>e�=��3x�'?�7������|�/`�I�vy�tVr�}���˿�N*�񆙥һ�%O7|1��\̖pnd�e��aoi��[��G)�x'߄���� �i�>XQ��:�(��%x:�{7Uٜ��i3̃�Hs9��L>�j݅ށ�X�~����������qa�b*cgs�+��*T�BR�K��G��Lf�t�6��y�h�ʯQ>�OE#=2�A��Mu$s�#���"�c�Tv5�O�`ʲ����)����tƬ�A	1�-��������~��&�[��*��\�bӆ5سc;:�aA��ܲ�f�U��;���������	�:C�tU~��D��?���gc||�����O<!�+/��3$�rI�K�a(C��K��c��]yp3+C�gr;HP�	�5�__��)�(�f�~��\!]�c!'%�V�������p��������vxX$j��j%+�V�~fa8IF�d�G���b&+�U6� �Kr@�-h��^V��Ϟ�o�YG�`?|�
�
*�RK) ��zn�7nP���#�b��<�'�ǔ���e,�\��t��L���+���(\@�3>S�gi������vai9c�B�r�5�I�f�,�^�
�D ��S��]rq]�����p��j]!�V�����"��Q�z��"��q����b�@T���֯Á����Lb�uسk�~^��7o����	������#:֑h7I��-*V�8д���rfb�	�4H�,\y�|��$B�b�t���=�R��b%_�i,����̠&�G�6@n��>Y*Ȭͨ���
)��4�=f�����1iQ�)G�V�ӵ���hzx˛ވO}���0���+.���o����wP?�V-�w��.GWG;����X�y��:\{N�<�����q_q�~��,��~h5����0>6�b.�p$ ���Ǉ;n~�ؓF��G��5X�y��C'e9*oy��aqf
kVu���#��p��s��_�UW]���I� �i�s�+^�O�sx��q��\s� �:�H�}�����?��� ������1�1tO� 
Ŋ��O=sW^s=����OVg�I���v�چ�ILO�j���AJw��%zA{G�x����ك~����i����&qׯ�G4����e"�ϫs/�Ikm>r�6m�?Ԇ�����F|�OcdbZ��\�"��<S���Z��N�:�o��(�B�y������][uVrYRB~��Q��p�Cr^{����"H�����+7�����B�2�2D�Y�p"bHb�� 
�k���'o{�}��o��Wh�^���?����K�{����fK��)�����
�T���Yd
TC�7 �ÕI��Lv-V �.s+��DTB��3�f�C�:u��橔E��ܝ����X.��38��9��Ym:d�E�v��Tj"V		�FbL��5~�ᡎ�^�R.[�J��H�V�yy�q���Y��5p�Q�]�q^nL�[g�������P�@�	�D�&�y��Rwq��AY0ǆsL���E���<���<��a�E����>Ҥ�2z:X;4 8�!w�QOON�;�V���I2}�%�s�ngYf���٧���r��$!�����A�3~��ϙQQ����� "RE���B ���{;9��sv�����w�w}�|��x�r��}�~��}��^�*��z�j̞3K�n�찵�,?���aDc	;v��^}���<�T�0�v�-8��1�����z�&��w�=��RѤ2²'�BuJ�r��7͵e�k#D�X�q7N���5�2$P70��:�y457`���z�!�hx��	�i i�/��3IT��P�w#�e���ȱ�*�S̨�����ͺ�yq �0F��	�ˤȔn\����䅰������p��kN�&�Y��+~���'��������;��f��99���N|ƴ�Zs<�T�岂��aOj�*d���e�U���,e 9�*#gE�=�ܐ	M�E��~OYE�~'B�N�a�����^��@ r����0��QkWaz6���F�F�΄I���M��93�����Q ׃��m�D��#Y���_�fν$�VaC���?�+���3s��)X@hxH�O=�8�X���N�����/Q�B�$e���P�hNA�9��2Ne�q4v֥��4˃E`
�Ζ�3�]��,D����V,T��N�aE�3Fy"��Xp$�`�\|��_���<��{�����KW���A��Ux��'M����YN�˗/����Chhi���kp�����I��^��K���I��������E?�TgU��������m�48�A$�y̞�?��C2�d���{��3'����3���W1������<t,X�cǏ�ˣ���C!���6����L[YQ�e�-E���-�DK�8R
MIƌ�f�d��56���������m����+��~*>��iӰ`�5	m�12<��Ml3���������)ۀ��*��Q]ߨ������ګ.�P_���Ν���v˚�A�\;䋱@c|�Q��݃P,�s�_�?�0ڻ����%��G���2�"�!�q�>��XӧN�ܻ���'�{>c�4��>�6e2����}��R��T� ��[��/-5� n�~�W.�@>>�R���?|�/��(T��ƥ�/vſN��� F�yE��Pw1JIp&�"��7��eW�p�	>�L�t���,�l�l.d�3(2f|Y���_|:���X�KP&&��G���Q���T����}���F$���O���R�N�Tq�S�&�RZ��Het,d� �s�'`9D�pR�d�:�pa�,)Q��7I]?��,B�ȓHt$7Aj�<.�`���|�Ę�EO4���v���#���C��I3f
&;�����S��&Cy�+~�S�?,"�Fu}i���E��e�/�E��f�	q\C=\t���n>'ٮ��ԑ�z���тf\G7���Y8|~9�2#���-t��(�mrsh��3k8��֟�C�l<�A���w(��H@U���C�(��@�ű#�PJ�h<���?�7��^��X�Q��QYꗤ��n���B�&�\o@0�Һ-9o<q�늿�=��>�n�5LwGGѫ���B�r����M^e�"�&b:�E8V��蔽z����%�dlv9�ҏ�땾F�Dͭ-x��w�n�z�^})�ʫ�֦wt��)�?g.�+J���m���O��<ɼ������PSW��G�(��څm۶���	K�]��G���H�e��H���h�8o�<�8}��f�-����C���D�p�-��眣������)m�7(�$����(� 0�,�r�h�Y��_f\ePI���((�N�X.�Y��׿�ۛ7��O�V_�T]�?X��p�Ca$Y,���3i*�^�kr����P��P�Ɛ"�/���#K�,X��T���l��nqVkL�{�)�,T�/��{��%<����g�N�VV��*�����X�d!܇];�J��}��
>���ή)�h4��Ջ�����<��3�n,?��Y�{�������-��a�qM��n�̙%�tǮ]h�&�<��.ÿ}�~���q�-���~Bk3���o��lj��W@[[&�M��;1��Yf��n��N��������d�p����:|m��i`I�2&`\C<� *j����}�^���&t����<��Y3�t�|����,�bph@������\KTKQ55EIYF�YT�6�G�����
���_&t������qFrx>W�d����O��C��]�C≬��J<��8�Ջ��%=n{,�Z[�UV(Ј-�}���{��G>*�IO���a���&���rn���X��>m�MXLq��G�
��3g&
_66�Z��_��C˧�|�o�?)�r�c�!���J�N���� F�*����Hfm�����E��M27K���G��,9i����F�8�<��	I���X��"qFF��@$���_�x�xF��t9���2����9g6Ot��͐�<Lzf�mo\�M0"*ȧ����a+�PQ�G:��k�5�%*Ӈ�t0�tIsU�]�rSC�`8�Y���E���	2�K4���Q��\}�F#߼�>l۵[�)������~�U��a+�����p�ܛŏ���x��\�T ���У��Δ�Ҹ��;��h�"K�B�1��� A��1}i%eQ�9{�`;w�D"�:"ǡ�?� 7����Uɤ�,��I�%��!%W�T������i^$>C:$ς�s�oH�ő��k��D���ey`����E��}5�c� a��Uک3���N�L��t��F��B�d�DxҌq��k�8�,W]�@|�,�X��:������h�����&�&UV��Z��Y��\S�P�
�.�m<|}���
X�p>V,� ��zS�u6���_�iӧ㉧�B۔�h�4��� �/���Ηw-�o��&�ܾ|��C�+W����;�w�~y6pr�1w�B��׽�{q�֬\�뮻NFTgN��Xf����)y����Ku8]E9��K�~�}�)�'8�Y\�l)Z����Q^Rb������p�"c��0�;L�f�XVQ�멵��!Bޗ�H��Ir�5�2ח������|�g?�	�{���"���?X��P�([�	�nl�|&��� ��X^RES�O���G�}Xxg�B	���~�Bk�2[�V�E�%g�ߒ�s�|�s����~�C���-[|.Z�Mƕ�]WS��>xG=�좧�=O�++��F��n��.����'��5��K.�C(�.���q}=�GFEd��Ƈ#���T&'����݈�Sf���L�_��x��<�T���r}&"�<�����Y��#+��Ec����_�/}o߮gaj�4V���,��WE�@_�I�Τ�QVV�=����eU��V�_�LG7~�ȣZ7��1�%n'J^�O�tk}��1��~Q	(� 5<F�p���u�Ƀi���:��	�5�(�%Q��32��k|J�<����q�k�s�0j[����|���Ee�7�F�(t�2���#8@T�(9�Nq+N��E[}6z�A3���d�J�N3N��T:����q�e�l����5D��|��0����;~�gR��b��_����"��T\��GS8q��#1����flù#��T:��Y6>�L��):6">7"z���,Ĥ���    IDAT	�)o����!�sN��Q�I&ϼ���<i�h���o���C����7#f�f��O�.��B�l�B2-%�)�,��Hb`�_�$+k����2c�3ڐ9��*�i\�*V*Jj+��^[Y��S�q��K��[o����w7)��ΗWa�g�{���A��H<+GG�ӏ�>ަ�?}�[�BGk,��h���.5���$:��7�d�n���a��*
�t΢�^E��f�{�drTI���Q~LY��'tp���$�*�+��RO���{L�@֨I!�U�K�����0��t�E�,��@�"�%?�SKEAކ���H���$�ʽ��,\	�g�317����(��b$��$���D>^+�c�y��9��<
�|v��!�F,^7\>�8.t9%���C�כ�?TA,�SŹ���9���ᕣ�S����Vn�M���K�tѹx��1�ߣ�7�+��
�����	�PVV��׭��IlK�[�n���ǧ���v�� _	����i�wt`㦷ĕa�M���u�-[��>�]K�1�m�_��`�P�g�`�<��]pх:�6��6P�ۯ��jT��੧�4k�� �fNmÊ󗫀�����E�a�UWa�%���VZ,�첂Og��ɣ�ⱅ�Q�/�sO���.z��Bئ���v�����cc7ݜ���T��J�xy��14�1�[�m���X��,8��u���Hp+*��o��ܗIJ5����*+�C���{��{l
�Ι;��}����8�����A�m�q���J���ÖϪ���"� v�.U�5��D�j�d_�?';�g�{Y6a4�����y����F(����j:�}�"��E���%Gٱhw�y�L������2�$���CM5hj�EuU��3�O+�?���2�iuv��ghH����ǟ���	�WJcufL�$I0�!{rBQ�ܰ��/H8�P�7·�}��q~�G,�T�� ��6��c���["����3�݆��&M���#�n\�m�ol�?}H�_�G
L�W6��A�Kfr)Zē�x��"U!�5���t��s�����=�8v<�)J�3&��ʖc^�ʑ=è#��ڎ[�l��y܏����db	�
NԹ���fP��'�Z��ۥ�se�H�-���禇gά��7@�ٿ��"*G;�c����Éτ��r��$O��8v�=������h��.�h{�NGd�lW�2����ual��XD���)	nj�ô)�D,���,�a$����Cغ�(R�� B�,����iu�<��#���B�fHY#�����)~��E�@�d�:�8�ʘ�b�b�'�~ds	��Dv�c�֦G"��9)�nnnU��C�jV��aL�<	_��.L�֊#bǶ�Ա_uՕ:��{{1��}�{��P�2	�@v�;�TM!�]0N���ع)Z���4V��YZVЉȨЖT,�|&!�f��a]qq�k�#F&s)fdD�"�k�9sq�W�o`G�����G��Ԭ`����v=D��U>�>����XaJ0��!ʲ�r�|���U�y8@����dl���$��}�F�Q���{b�tӉ4��$I�u����b��{񋜙,qO�[�q^:���E�F8���|ߩ�A�=��|2<����[B4%�CUY9�����RqCR��S�����hS�<y*Z�[�a�)�����K<$��rV����k�9��Ϟ��(�,^�5_�g�y�C�&C+���W_�#G����	�['��[`���u-]�LJ�}���n��q��o4�nW�mWO6n�d�fD��9̜=KΖt��[,S�gN��77�Gh��Ƙm��Ux�����TZ�S��@^t񅂥7�{Cv���`�3�>�_}J|nq�(��a!�?K�]���M��׏�*��H	n�,L�`;;�sC��,*��Y���c�7����ԩy��ₙ5�@)�"	�D\�τ���u G3�x��I�r���y}";6ͮ�e�W���Ҋ`o!&E$��m��}q��8�-��/~����aώ�RaqoeA0k�d47���`�xv$�����'���XL#��X��$������?ކW^}M�9���k��*��D4b�mȵ`��͆�����1M�Pa!wŕ���s������.K�K5T�'O����0��kcT1�pu�&3f�Yt�� ��`��s��Q��-�&�aC6�ܙ3�w���ny�8��s�k>E��.������?��c�A����E��'�0�xkkk�w�P1�C�Rlvk�gN��o��J\{�mh�0?}�g��@0`xOUe�(�e"�XWm�X�O�$���e
Y�Dw?±$f�[�kn�	O<�[�wu!��$W����
�B#A?��$�l�9I��d�����%�
=L
���Q|�{Q\��
�}�Q�+���&���o���9�6c����'-T�wśéo�%m����T�-rO(^��S]8�ދt���}2�NԐ6S�0<N��aG4�c������O���k>ɂ���Ӗ��7߀�'�E~���p���D��3/l�G;����͏��<%�����Թ��j��+�Q�D�,��@�����K�b`_نkTB3��HF����|�D|Բ�f�c2:�A�»�1҇��~S��]23���+.ǒ��0<Ч>���H�2��A�[��}C�Q&I��{���r��{�Ҁ�\�9�`���d=%iAI�`�w&��dԻ1�#_%Ә+��������@�"n�
�$	���.�hi����]�]��`ۮ��FÄ���8��a|p\^x���"��>`̽�����F<��0j#{֨�┸��1�zE0h����
h,�c� "e�<�IvNm�"$Z>0�����ɥ"��P����D������t���.�X�ꬱ�:q,_7"BT�8]X�r�.^�͉�إs#g��n�zL�5k׮���(�~�qAd�ND��u��1T��w����e��ѥ�\����m��p�|tu�+�h��=��`�9�c��e<�O��o���̵'�7y+�0�����={�s�yOl����l��c'���%�4w�<�,���ǥ !���F� 9j$.^t.>��C����G�`L��s��w }����i^@ei �^u�d��O�D��2�dq�h���T�U��]4NT��B���@@&fB�,�8�e���8Zd����~��~�Il|s�Y7�u�[���1M#�ʡ@$�cN�=��/k���S��Pcd�)�V#K�/߄뗖�Pj��>��$�v�p�������2c��r��x�d���:�k�Ʒ4����xX( ��qu��q����Ө�j���غm;�|�鳼ퟹ,��k���+K�FM�5
~���S�����[q������{��ɓ�g�kT�"vbK�F�T.�_�E$׸Ҁs���U(`�9��׿���ؽw����y�*u�8�`�L"5�*Q\^;�TY�3�D�Î�}�k����#�?aƃ��h�IUUV��p`�Vj�� �/�?�fxdhH<$��Xu)��'����~B�s���!���5x�jb���.5=lВ��
��/��܅�qͧnă?�dy"��C(	�i-�ژ��{�^�R�&���gpU��2�,pD���j ~���^x����J��s�=���z�%��z���d �O�F�������77>������������͡X������#iwI��ENGs8�H��>d�d{�xY�J�~�b�a�8�����s慞��4-b@V\���iS��S�ȶ8X���%ԡ��'��w�� ;�FŸ)�?ѴcqrWX��չ����$e��Ό�
i����-�f�|�r:��G�6�h�@WZ�o,T��B%�`��RQ$ҮQ�0�k9� Z���!Y>��ǣ�ƌ�mX�h!b����w`L����W���@uU=�ܼ�v��GP�8�@	6����BŮN���|�M��SV��D$]�R6����y�#G�i�!���Ò�G�O���mL��Y��mq���Hc+�=irt����a����Xx��.x(���̘�8ڋ[6�A:hi���]�."Y� ���D@��-�<$�G��x,��2�A`�����/��m�a���$M�+`6Fv��B%�cg�G�*v�H����hH��bBˎ߬ �]�
�#Y�ח�Y3Tt�r��" .]����aͅ����z4������'O��q��'���3�Fnms�}�U�5
(J�-��b�GMπ� ��^r�
��g:�n�R�(�GN	͞8*�Ke(�H�)��+�9�h�vy(��͍���թ�\#n�,��/<�����-Ċ+0s�4�����yr�5c�4,?�|<��38����y��i��q�?v�$z����٩uȑ�'XP/�7-��4�<u�F\[D��-;ӧ�"PYVyM+�$�PaA�g��PSK���I"c>g�K��s�?���� �}'i1,AUM�?�8S��)��H�L��a�����ds_D�5��v69$��b�~����q��KⳚ�K6��,�(��}��*���3�|�+_�OxPq�����X|L�JI��\.��+ΐ�$;�YN���u�����׿��8�~?��?t����#~����4e"Sn���:��c'a���O����?���Б�VQf:}�K6���+~	U�a�*)��B�N7�̙�O�N����x}��&�(9ɢ2�4�;�je���xj��x?�sn����o!�����1q��� %�=��:��Il��.�������~�k�`E����S��F�$��y����o��$\=e�Tt������s,���[p����c*��5R�~E���=Ʉ3�H<�<G�N�+�B'�|��d���ԩ h�&�@	~$Ld;��͉D֦ N�?A� X	ȯ�؇�%���	Ձ������E�r�T��?��N8�X˺KrJO�����هށa��4�*HJ���i%'�Fz�y���-����:
71r�	�&�������ME��q�K���ו�ؙ8{�E�:Ўpڃ�ƩT4``4����ql漼��H����,T�a"�/7�_up�1���0�\J�J*:�_
��k�*E'�tF� IM�[��bL"%>�+�-Es�8;L3�1T��JM�õ�UU=k�<�^�onz�~�o��>jƵ����|�� Ib��Fi�.�q|m:Q�ׂ�t���\J���3��n#�@�v&�M��TJ�y8�����.��c���O?���Q8<>E�s�\�3c>�$���Y��=Y��;F��
3F�Z^�<�| �1XV�̄6�p���\���Q�����<:2�])�����yp����n���TZ_n���R�(��6��;D>2r�J3����*�O�bFo�yL�e��y���_��-ǃ?}@?��.����v����pɚ58g�|<��c�n�����b:o�Ly�+Qܜb�1�5DβjV���-Y��o������T�����:\~啸�����݃ݻwkCWW��'O��ޓ��3g�g���N����E�۰q���9���g�Ξ5G����+��R��S'k�3D�)�mm�p�����?��e�ƍV��C%�6���pp䪜O3�3�	�"����� �.���\:c��=t]6�NRyks�rg�J�-�'y?������z7������(��"�u�ơ��T��x�X
�,���PbJ�JJ�9�4\�=��Qv���A���~��{,V��r�(^��	,��,��XG�p��D��3eԓ�?Y�p���0N���6�_��qIЯQ8GE4�R&�3�"2K>�A��_ҝ�������~�a�ۿ����Q!�,0��cT���ؘp��B�.��|�sw�~\^z�u<����4���2D�.iɼ\c�؎�<�7�����{�*�;�;��S��ѣǵ/������Z2#Ӕ�J��5<&�t�eQ�����˯
1d!̑�G�aK�e���F�ET"e��.<+.�X�Y���O>�g��
ݥIO&8E0"�G,T�ܫJ|j�X���h��yXq�J�W?���%'g�%+�ҀF8�* c�8��p��q�WTJ�L%��C�x�����ȝ��ӡ�E�ɏ�'ԻlG(��h,��15�-L��J��
l
�g"���j������G�k���Qa�20���X��X��9�qO�=����1�*�z��d�1 řG�u�b�TW������zL�҆	Z���Ь���T2"�ݍ7݂3]����NtDp�D?�RN�4M��W�H���4B3��
f;6:,H��o;^e��A�C2P�#�LD�ʟ\����j���+��a<�yhL@5��<X�,����e�Ƃ���Y>��Kif� IƔ�q��l�䦱huMM���[�i�;8p�86��J*jP�،u�� �Ξ���ϊ����Ŀa�UDS
Ƌ��h��p�57���g��� /)��i����Ѳ��)!N�"PP&[prP���>��츉���䃧M�A�Ҽ6�b����DвMB.+G^*���C�9��`Ӄ��}txhp3%<O�I���Fgfe߄W=)T�8�&��?����������K�5X��}jtF�}vc�2�_�E��rru0	�3O���d@FW�<|.���t���������L<�,\���+Eկ��R,?~�sζ{�.M�0����{4�k|���h�͇-�T'�b���X��duNg_���J�
QY�l9>������=g����k=q�P���Z[[��G�H��pf̘%��U���u�:y
��+�g�n%�������_��m��3ɺt�ͧ�p����"�I�lJ����
���s'G(
C	g���K�`j��I�uu5(-��ʋH��!>�p!�S,����cغ�#�ܳC�Y��Z,`9�
��#M �H#Ʊ�Z'*��Y&��mq�#%� ���P!q��(I�I�%����� ���4\JT�>c�"���T1:�K��%n[K�]��o�	�N�� �L0�AV�R|�������JT8h���I<~�D�:uu������?�(���Qz�ﷸd��g��&���g�P��ӧ0�|I�9V�?�F��&���	����C>�X׫}��\�l>��ߏ��jL�>;�n3�`6�AYmD*k\d���Ϧ��	�ܙ3w�
.����׬�T�5*,��B����=���:����}����࿯���h�<������U���ô<og�T��L=+�=Q�b������G��/�fԘv��V^r�bOj�+���@z���~�诱��ayq���1(Qc��$y��<YܲH��=7�,��q����1�1,V�R��H������ÖS>30�������Ŋ	6�?�Y��i�'��ߐ�{K2v�T?�}C���'�0�:�c1�;FO�q;�Kc���|)ʃDRXyɅ����8v��z�	� 4ҏ��vx=vyIP�C�c���y��dq�+�dރ��6���$���yr �b��j�#�����.XpV�P����PȐ?C&1
G!���Z�"����Tu^T�Y���̰�1xƷ
�%�[��H�t�e�18Ѝ��n}~n.��k4_%�.��ޗ\�
���9q
���DiU�5���9?�Mo���
/(*��R�m��pxغ���ч<CXǥt�����r�0#����� �,n*^&�M���(�GBp0񖪞B^��
A��E�;!FF2m8(�^�[]KJ?sR�D̞9�U�b����w�c�0:�]{wa��6\q�e"�r�9v�0^y�US֏����]�ķ`����ٗP�|^�~$�a|��1�"ac�N�����e�u֛��2�GQ=B�Xc'B���4sY\�j5.Y�R�K��mz����o	�Y��<\�j5~��/p�����>7	J�"J�"��d��%��k=3)9��FT��z{�(CCC�)֝��V��bqE����T�����<���Z9��FU����a�C���ScCm��S '�%�a��R �Μ�;k    IDAT^;�eM��\�a��cQ���`� ��ynN)��?�cq+G�lZ��y�x��r�e�]��M����&R)E�G������?�P�k��
ؔ�)����0�
�霺O*�l���Q�)�C���!r?,�|�f-cBU�P
�1�_��+�<?�P�aC�?�5��{��a�M�*Ә��z#ϑ��/�@�DB�g|f�3F#cz?<�8Na��kA�!�{�:�;���C���f���W⿑ߑ��7D"�y���5ؔ%�p���A$���F��3�g%�l&X��CS[_����A���o�G%�j�*@���h"��P߈Y�g���
	Km)4�♱U����%�s:|s�}�N睻X랟��	��.�"Q]o�=��Ņ_��!C>��c�Ż
�F0w�9���>�����~&��3��A�!r�JJ�z.GBػg��z[!^QkK#���2��x�L5�~��FG�4�S�L��[���-�9�T3)=����D�r$������$��q�������'%����5o���к65��x�^�D�;)O��൥�Z����������'�>Q'�7�ʟ�L��;�<0�^,�X�B%U�b$�U�w�����	7	
�E�I/��߉�St���.`ْ��,B�Mu���`w�qxQ�R��~�8��%��o��9����#����ɮA�;ډ����0ř��5�4���fl�_n���WD��y�׉;��S�ņ��.�h��lr{Z����R6o;s��1�X�@��pf��ǑM�4sg�r�uWˎ?66���^ɓK������X��X�h	�͜�_z���Ɏ^�46���o��6"|HXu����,T��+��c������	"a$�K�h����n�~�W8�L�5�R�;��ꦛnQo˖we���ܢY.G�Z�fM���Ň��"���4�al@�t�gp�����Bۤ�X�j��"F���&��.�w�ޅ�^zI��O�ӖQ_�h6�ǎ��0c��z�m���X��zlظ3���-��,�x"��X%�%2�r�<���+�];1��v�T�P��4kyr��ټ��hvk���1˸��m�C-<~��W_�+.�TQ�<T�Q3��_���G�鯹�J\t�*<��鷺��I�4�������uD��(T�1��fφ\L�?]H��B$�J �viB��^ul<X�FB��DO �c!��C��]#�f�|��\��Ҭ����Ź=g�,$����V�x:-՗<r�8V���T�S
�Q�py*�:!ǂ�4�-��j�@��%���2I(Ϭ3���t�)�E+���n�������IH�I�u:�暅]����*q�Ɍ\���2�	�s -@ҿh%��z���Y�4c��b�����Dԑ�����ݩ`c��0K�Rh=/�@���5ry�}.3
MfL����M֐�?��q����'ǋTװx��T8Q��t!�A!;i�e�"�NIZ��N6^7B��(-)��?y���9��)-ԏ?�b�7"o��l!Ϣ�{�������I�4FBX���W�٬��(rS<n�^�����My/�eez��Y��Y4(�9{$�M�4��D쭑,	�w��y�áQ����I!��<)��PQ�b�Rz6g�R'��؍�e�'���{� )�����ڥ�9�+/<���y}6<��3x�Ģ�>̚5�D��������q)�������y�a�#
��7�S6I���<~��8r���Sv������i����a�����ϖ�k���w�u_~|�B��
�o"*,Tz���1�u_O:R2��H$��^z�!�HHB&�lz��"�=s'�Fb�~g��e����2�	x���5���1y6�v'�n���l��!I����,�7P��_i-:��p�tb&O���2��gc�3ID��h��|+��+b7j��ac���D24E�#��"�����b|�8�#æk$G�
�#��(���(�́J�H�M�4��˜S�켅�;{£����F��t��d��:,:w9j�e���֭�`��G��ME�&�{bTQ����V�d�y���X�A�D�$_rH��4/ͧ���-�;W�y��~��:s�3��y�&o��i��ʫ��b��k!�-�Ӧ͐���x]D<�7����m���Up#`�HO}].[���#$�n�GV�J�G�D�#���M7�(7R��N�9����5�����������B,�m\��(--Goo�
.���L�ys0�e:��������i+h�*Tx@h?�FH��ˋ'k�}xP�&rU�9��4{���q���#��5�t�,9o1�y�=lݱU#��W\���m;�ˡ���K�
=� J���DEy�) ���4�RDG�T�q�s3
��h�Hc��m��!sg�B���U���;���$
��UTK�7���"E���m�g�ad�,>���B<��� �Z���&���L
G$����E�<�*�`��Pќ���>��/�0JbY(��O���DM}��c�-x ����¢���ڰE�%o�*�X��F�6#�5���c0�_�m%Q���M1NS>�)t,��b� ׍�?O��H��o��l�ap�e�F�W���uZ�å��nD���q��8Y�[���n�/Q�fx,v�����b�-R��Q��^DH�,r#X�P�B�(�2X��9N���U*��
�ޚ�#�c4�!L��of��L��F�Du�s2��:�b��\�D媫j�,�*��������N���Y�
��s�}y� tdĨ����epZ��T�����
q-�@��z���)�	��&~��gF �}���c�<I*jj1��s\���L�ʂ�
ǖB��5#Dq3�;�h��9����>ZB S��.Ǫ�ᮻnDǩ3x�7O�Kh��Eʡ#j�}�^��p�=��{=|���d&��T�'����ƛn�QH��ￋ��*����_�(�@��G�N��\�\�l�X��D�#Z�$�gz�W����O���ʉ���P쟒9�u)[I0�g8WN����Q*�4X�ӏ$Ʃ���u� ܠ[f��sf���cG��׭�������ǌ�s0q�D�ڵooވ��5�U*�Cg�T�WI�"�"�;v�g̅�W�H�3_�60�sP]	 ��8'tc-�AI⢿���.�0=Z/�_��ƐKD�g��T�pxH3o4�#�3f9
d���ӫS����hD<&�r�#C�n�i�����Cpko�^gϜ���a�[�AFK�v�G4��ܥ硢���߈(�5�DJ�
k���)	�$ԟp�$O)`�U1�*����VLi�����m4Lz�C�M���o�]	�<�6��	�M����V�,���>s/��
�C#r-���B��-��I�HX��ڊ믻͍ڈ^}�e�U�*Vxh� �@~�ԩS��f�v�d�L~UQE����[��p�s뭷j��A���O+o���N�T�p=����ظ�-��
⚠������,h��.TT8Ѓ�R�H�΃V�G��n�7��S'O
�^�j�^���&L����4�?�ف-[�()����L6
����4��~�ͺ!��H*��tv�#�3���Ș�+75�-U������i���c���t��zfx���º���\^�6GA��Tu�H�$�e�ɋDR���nY��+�t`�tIw/��
TQH�"��R����DEbF<�8f�� �@.J")"&yP�i�'	�Q��_C�	D}
��lIhϓ��j�邧�\�)9��G�f��>�/�J9�ʲ�I��)��x�̵�CV]z1.���\K�%c.f;+��"��
��gj�8V�ę�Gf� �.
j��X����VN�"r���0����?8����l�ܝQo�wn�޽{,/�y˗J�1a$
���~���	bG9��,p��9�	ˤ������X�3]��S�c��ɨ��P��\��s��<G?\J��\��N�Kԍ��g�|�����k�ZД��?�6l��爫*���ϭ5¢_��<�G9v�>��b=n��L�8Q�|:uSIĵ��'�v�	%�B�!�|�Y� <:��h4���u7Z&NT�E�Qwʒ��P���C/�%�DPYL	Aa�X[�{_(�x1�(���R|�w����=���p�5W+5�E��o㣭;�_�+=������~���U��~���\t�b;~=�S̚5C�(CN��o���)��C���E�gk<E�B6�̘��B@yr�{BM�[���_=y#gw���?��g��������+�ʮ�{�J�6�Gsf��?���� L���PNڅ���'QS��M�_�����xM����
��(��D$���W�j��0���n�N:����U	E��� � ��c�����`��s�9�ʚ/C�R�Q�aDC��%#�e`�:�>˫t%+�A'�H�.*T�65�"4:���>�$̐�X�0��X%���:�L�Ҡmixh@>*��ɦ�X�j%���J��(/
��58�م��v��������KV������B��P ���C��B��X�ɑ��[@wBC5���DR*I��¸��j�t�7�'�-��iV������r,�j�u��E"�tvw��·���_P�.��2|���l�6��v�lhg��X˖,���ܢ�h���x���+}BK��><ى���*dj�j5�x���W�P^U���nu S�L�uݱc^}�Uױ�⨢����կL���bڴi*z*�*��?�_>��Fmc8$�g7N����TΧ����e#A�k��Y Re�3m�i�nch��.+J���m���аE�=[�X�vv��L�]�����
��[�=�L��lT��r�vZ*"�}2�(��G������dLq,b�H�F.k�)��(�m�!�=&U�n\Bc���-�]�L�3�(l�������/Ҹi�
����!�25��	���}b>�v�<�7mz[���i�޲H��W�4�H����� NB�';d�W�/���x���F� ;d:x��hy�`!�k�A���["�D�,�d�b��u���J�`�aj��đ&g��Q��|�^���S�;x�.� X6[<�����T��C746��	�1c�,�ص�� &Mn񙟃�!���d����c�M0�)��[+�pdSY]�)Sg(��xK�x!���ڋ+˃��������I��CcW��ļ0F@L�1����:a"�8����	�IQn�p�ay%|��A�[ �-�6��oŒ�KUX2c�ghXdn=��=�z�\7�2�Vh�Ft��k��ɪ����E1u�t}N��on2��4��C-�
���9g�D~_"G�Đ�yM�:����o��Mo���`.��Khi���v`�GJ�}�W����m=��=��������O?����>�9q���:���X��2����w/>/�9�.�9;~��3�y�$����Ļ�A�	a&���=�qڅ�8��]S˿��?����Z���ן�P�vb��{`�3���9{iY2��p8���a�K�(H�B"��P�
�����;�����󗢶�]��V
��'NPP����)�		 	���S̈́��TTUax8
��󖜏�Cx��7��c�y+1g��17��\<:��p/{ڑ��P����J��^x�e�V�I~��6uo���f������P����z���s`��El��f�J���iİ4J�8�,+	���Dlk��j�1�u�ȏ�t	����"$�d��XTp0+��3�`�9��+�Z��� Ln��2�Ӗn��q�,�q�9[�[��\~�GV��HH>67�p�B�~������>�6�D,�M��w~F�֭[��Y��l���+��&������0k�*b3��fNɰq�$'�]7J�͙�k��FE^��v<��Ә7w�~��p4"�ޑ#G��ɍ�Ғ���B�#B|��XPp~�u��K�,;�O}�S���N��_D4S�@�=M��k������/���^�w���%�$q4�£�<T��T�wC�sX�p��1��;�B���0�17z��xV��q �Wq���\��rHjV�.���L��<��7a�鳑 �&yT�h��j��!���?��d]vv>_=���4\�Y�^�9�gഞ!P���u����lT�։���D9�	�4H!��EdN#5��(|���e��XW����-�_�x&�^Q��󪰧���%KT�Ҋ���`?܁��mm�D{�E
��;L�!��,r8�"M����?�W>��rID���[�T\;��2�⬱�Ak�FI�����q}��G.OEY ����TW��������/��Z�X��q�2��qR#u�S���g�s�1��W]�{��9�n?����Ru�uY@�x��l�8НU����/Y�_$s1~b������G��o���M�����Tl�X�h�KM������.0Ä��X{�M��+�������ѕ׷:`�fmmƱ�A�*�R��J��ż2��H`A��o|����O~��G���_�G��e�D~�ǫ:Q;��uO�ڲ���_��_)��=����c�F�d�OT0�,��`�g2�#+ͱ4���
6\s�U�>{�z�Y>qL���^�P;��`Ãh���wӛ����crtw�lx�7�a��=���/c��f<��+��ڵ�c����4�b�B1ʷ��s!*��śJes*й���!��8l��pd�:��W�Ë���m�D�_�B�(��)����JJ��8*��U����Z.�p_;Nލ��(q�PS�EkC-*ʃ��X�J�h?Q�qHdq���;ؽw����#���r#>�sPSS���A���������W^G��Ǵ9K���a,J>
	gIDG��}Ý'��8�*�I|��=A�V��WZ�B%�L v{�>'�K��:��X�B���C����E�:(8�K��3��u�0_ey)j��e���խ���-v;\�|��rS昂�]�$�;zM�0�r̘;/��2B���r�T�{��I�������$V����q�2������\|��؈�)�����1<8"V?����>��/��y�Z�Z�VT$"n~g�� ����ŗ��!)-�(�neՈ��QE��H��뀤z�ĉ������ѣ2kil�ܹsՙ��1�ӣ��3�yV���Z��bǶ�شn���JIfى�r=m޼Y���E�8ɼ�/��3g*���	�ĳ/�V����lvm�DT��5g9.�6v�)���q�H�ͬ��x�p�e�-yP\#�HXELIY�Yc.�9�#2��qdB��VXc����@VMa�Mt�a��b��I�����z��t|��p�-��9�1ȳ�r�-��~�����~�ocx4gQ�PQ~"�\���y�H���×#DFНU�=���粝-TIY�Ke�a(m'��a��-�K�I��ݥ�R��pH�
	���Hy��wq��sM�$��`M��$�	f���`r���'��%�Za�ܣY�"�KP�;:ɯق�X*N�*V$ز2>*TT��8)+�3�ON4�fj/*~8�(���ݝ�b��Ÿ�[���7��{4�.���k*�{��]D£*x�1}G8�N^�_ȥ�?-���w$������2K�=�1)��������ɦ2�o^�G�8���"1��_}��_����h?yJ<��s�8�n�&M@E�R^W|?,��� �8�����]�Xr�r|���~���gP�>2<�2>�vrI��`�yz�gs�#u�4��<GF�F��T?��c8p�(~��G�V�bQ���:G��F���^�K�|.���6R5��٭�{8��[oFc�x����L�"X�R�G��5UHI"��c����0�Ey��p�,�����������jW�\�ŋ��<(Ė�BGG^u�Bc
�$R���Ob�ޝ��gnǢ����o�þ}{p�e��l�R�;$$s�������q�g�t��ʛ��;\�9+���Q����
gf�cjC�߿�O_z�ϦP���S�Yz]�UL�8�Ew�0��C"M�����B��>u��.*�T��Ǟ�    IDAT��"9�<��4�ر2�"R���[om�����3�	�H�7c�t��:��0m�|\z�<���ў�p+�:y6�#LofǕG>���@z�C��`K���N�<�n�]���z���(J��h���c*TJ|N���
VZכ�X*VW�N�f���OFy]M��M�x��C�]K��x��3yOpl�)"|݆M8�~�\��F���E���[�%U)զ�7�/Ƒ���?FT�9��ga0q�x��p>
����&���!޻s���;�.����k���$+횚*&��nX�^�,z\n<������`�*��0]'lvd8?��t�%��R]U�;n���-*�w��qY�/Z�k֬�z���������_{�dg�����OH��.�<^c�Xh��;q�\sݵ*�����Iw����s���[��~,"����ZB�H��ъ��y:�ЈPv���ˎ�����\W,@
}~Y�E�3��|m��c���o�pVmP��Rt���"⤟M"�� ���z\�f�\�:z��h�Y�T��W�h	�캭��(��k{t�ga�E���lb������E:eҤ��K(�L��1a"�Sr����<�3h�|������G�|�#c�e� ����5�N�,y�(�KaUm--Z�Ey��>�HR��N�DOP䋰0f�����k+����x>s��(��Fg]>��*1pҐǕ�LT���I卓U�&�9r�a,�����M��<|o|޸�������#��X�����b<��S�loW�q2j�H��&OhEee ^FI����Iɽ����GN�DWw/Z'M���7_Ŗ�?�˯����֚�
�6�Cc]���Ǵ~��"jXUS�u}���F����V̜3�������|=���TD��IQ]^�A����3�kF�D
�=����:��C��l�*�8�>�l�'N��)m�ݎ�hOa�/}UX�����R& �^�u�w1��;��}���B!�=.}����ȃ$�'�-���(�4R�;w�ƙ�n8J�����r���o�CGg�P=�P,T&45`֔6�UUH���E�x���
=�B�ۻ��;��.Z�[?{����dg�2Ѹo1���̱2�a$"&�EO6���z2�3_Z�K'�D8<�
|I�ϛv���d2U�8/)���%K�o	\>w$�G��V��}PE�ׯY�d��G
�l�}Zc�7����<
rT�t�|�歼��.M\e�%2mH]�O*�T���ݏ��c��(�9�u[�d�b,X8}����&��Ё�`/*����Ҭ;B��X��#�����e5���=�';�.����K�O�qR@!���`�
��@lH���2�
�k����PV� ��\R2v��c�O6E6Ai�*T��G��"�1�Y�`6�bw�dYjܵ�x��M�9o"�Y;���8-�+}������,�z]x�j4O���^���?U՚�6�O�MN�	Q�g�t�B|�N�V�
�ڲ�I?u{�l�j�������� u����
���⩧��/�)J�*�!�"��x���7�o�b,yt�mS6�&߇�hvN<	}�{��E���5�T��(�1�? �#�qM�*"֭[��bF?�ػk7^}��_B��]$�UB���.6����u���w��x��M��
zn���>>�x��'�@5N�⛰8���������|'�yy��3:��V�:��H�?;vC^MRj�ob<:[���ῂ��J�;Bg`�t�U�d���b�Jlyk#��iX�����C��_JH�'#f�S�_gx��w��[�TS`�f���Y��}"��o?t<.H�#����2u\�3������7���_�^�	�;�`��6K���"ɓ�jJ���+)�ܹ���H����Zj��<�	ڸ������H8�xOMc`��YTE)�?�C�G�$��	Z��
�U.*p��ɚ�U�W�ǂܿ��b�C���٭ŪCE�i�fϜ�;o�?�������_�WSm5����m�!���BFDz�'�,y��	"PR�H,�����+�b���^�x�����1e2�+	L���C�J�%���i�,FF��{�0�Gq������oW�?�����0��E�D8�X���Ь��M��1
.�����	���;���/��mۑ�f�7��sB+�+���yFqt�J��>�|n'O��}k׾����W��5q,��㇐�uڄU��itJS���MsN6�|�����L)x{�W�1��ÿ�%F��Z�e�=c�Ҙi Z^���@/������7TW�}���Ƕ=0�����O��_=���D���땑G�Bvi����cw!����%њ���h�aύ"��{���`���������XmMM���ȥ�)G.��>qr�P4�2M�����
4:��j9���)�gz�AU�3�����uMm���s߽�ϧP9xf�{͵NoUY2���H
=#yH&j� �Q�E����m?G6�R?g�y4��Mχ9�gJn&%�������gT!��=)!�Ɔ�kh���V`���x�W�9AY]+�_u%����&���QȤ�@�i�w�@!5�LN�7�c
��[Z+b.%��V�r>-�f�P���\'D�0�
Bv�ȯ��Q�0�I�\��>[���e XEE�B�C*5�D�������RW%�s����ǟ�h1��O����!��� ͱ�*TX����CTP8���4��q�4����#���J{W\v)Z[���SO��$d�N�~�<k�[+^G2<�9���*b�ӎ���pT|�NjӵT0<����ҫY�1�'ƃ�X]�"�|/Ü9s���&�,N9�g��H%����$��̪�������|G���x��+0{�L�?��C|�}����{��Y�i��)s�9���Nz!	)���E�7Ad��]�]]PW��节�.M�� ��2�d2}�̜:����~�7D>�+��z���ₐ�3���>��w�pDj*r��	X��F4��7;<��tQ�EI�O$��BR8�'�&gA�0=v��ЄBrh3������B�pW1�{A4�\�P��p藍����'�H�"E*����")����57������W_�@OP4E
�sX`��d��UX_�ݡ���TˍT(���0�E$Wx���fK�Xu����nF#���R��F�I���}A�T��W��)^X,��+&Q-�����H^%��0*��E��r��UF�,Čq�}�"<��J*H���i��+���}�?��:����*0�]�ֽx2��o*���uH�FD��I��86��Z��BԔ+U���2Z��Ә�e�a'a,2YJ�K�����Č)%<w���ذ~-n'j�¨
��`�L$b�
$eT	�܇�����[���:9N�(��߅K����#���{T(�ٚ9k:�S�^Cbd�}��K�W�l����p��-���x���8��c1e��v���%S1L�<�gM�9�5,N�4k΃X���?пipd��1|����}=���z[��ĶV,�5a�K��@o��'6��O���$xV��W�x"�7�^��0�'ߛ�}��M�<'M����^�<�����y5�ܣ�gq�^��&L�9-���{�Z��2ur;/8Lc8���7�,��4Lgk�{��p�hiiCC�xlٽ�`5������v<�rD]KD#s��cD��c/ZN��9�T|0�(��ܥ�3gN|㨅�V͙7u�y�đ����ʖ�PwgGU����u;v���~,Ur.vx�iz�(�|px����|�<����Ԗ������������cO�-No�Y��T�s.���;8�B�P*��l虓�Be��m(����q��5�cN�����W����TVJ�1�hl"+�z$�"LR��<u����{�κ���	3�o�h�ȥ��Ɔ��C����Q��ɔ6�>J͂�Ҍ�J�7A5�X��%P�#p�P�F��ӣ�E��l=��B� "��!N����֢�Qnش>�Ҫ�+�^rTJ$Iʪ�B��봍�(�|2����k$W\|�24���?� ��Y۪[�U�8����s5�MA��bx��#�Q�bJ;�#�,	���FG�tH�C*;�i�钛,G&�n���/�1�3�<S�SO=%Άf�Ec��Z��ư���6�"C⬠���:j�7���#�zX�s�r��Doo�����j��~2�&G�"}!�N)���Q�CDf(:�¡��I���phâ�GX,XXH�(��Y��$���@��!�U�*�B� �M���B���$;����� �n��4�ơ��FV��E><(��z����Dk�m�ϡ���ʂH��$?�S�%�*1yBN:n9�~c�4z	qI鲝ll;�Z�pѝ�����Rq�|&���YJ$�R��p;��TWV�ҍ��8�|����FOh�׌%RR;1�����,J��ĊǐTB�"���H'�M#�������ON�e�ƙ��p�6$/�ƲM&�QD�3�y�����)8 ��kP#Q����0�Bj<�9�27T�*^�G�I�|~���m!��=尼
�+��dۅHe-��ը����K��|9�,r��	Sq�����9�w�ø�&���3	�:Ql�U�&.�}��Ի�G�³��}zq�1ǡc_��)�fϘ���͑��\@�rcz�Ee��HUX{:��[�;vtbB�̙���o7bhh�P�s��}`�T�C�H&2_���疹\D�������3Q�Ѐ����ˮ�]�ދ��[�ʪ̜ގ���@��h��=���2�}⽣g׮��0}�l�O��'�y;�f�r�w$�;g�̘�a�C�}�p���{��6OQ��˃ه�ǖ�]U֢��w��#���z`�q�Q`�O���	-HЖ��� f|�I`�t��#�<m��MS'��_����wX�u�
�WQ}�/e���e��q�ȁs�F{wNh�z�����O�:y^S�Ϻ��������ݍ����~�Ué�əb���F��|O@~B����NK�����ˣ7^������{�o�����;R��W :BDe}�#�'S�p�z(gR�ܳ{�o�X|^W�L��<n�?WFB����=-�Mضm�HS��=^�2�#���4��EcH��I�?R �U8�c��#o��β�L�+l�6���(�1�r	8�dIi��D� 2y�8��`\��(D��Vmm%1�����Q&M.#�W���q��T�;���N���h�Í���Rnth@ͩ4�a��ߏ��Zy��ڳOҴ-;v㤓O��i����O��p#�AB�uv,J�q7��f���d�#�����Ȕ$t�B������Y��5ˌ�PD�4�_�w��a/�&��:��P9�v_�^Vf�7&�AQ2Uc�E�?���(e@5�@�i0��Fi�И�ˢL#3U_�H_�)3�1+�#{���C� >n��'�Q���"��v�r�,���#i�6J�)wfwLO���z�?����Hy.<4EB���V�h���&�O�:h��b!+�A��i���M� �����ɓ�_캸N2)L�4I�ʺ5� =��"��%�?������u(5%��H!��Ʋ����mPEv��鄔hDKi8'���'���Q��+���Р,�B���!�4p3zQ���Fd�m�S�X�b�Z8�7�A�M�2�/�uK$��W�o~�Ѩq6�Ц`(G��F#�̮=v�S?3�ͫ�f����0�j�sq��[�<>kr��Q�&"�.EQ��9�TwWSP�A��D��#i��#�@D�z?'L���A��x2����2v,��c٢#qɧ.�]?�!:���该�ȥ
�1i\+����C����w��~�s�Ke��oa��y�Ɠ8���q����s��e�3sFG��P��۷�c�Nn��y�\r����3N�����m�&���m2fΙ�o��m����{Ι��!�:��׾�猶�;Y`p4|��c��k�X�[p8v�ݏN9>�3���D�jp��c0���tL��]��I�
��t6�1ߜ�S1v��s,�[o���+Vb,S���k��E�?gF��5m2b#��Qe,6"o/�5���j͙s`8�AMC�����q���*T�U�peȇʠ�w�>�R�Y!�|>kj�i��}!L�6I*�၇��{�!�)poʤ��%_�[�;��Lr 7g��	?����޼��'����{eoٷz�k3�l�r��g˞�t��/���^G,TJ��Cӛko<�Ƌ����Q��uG�͞ʖ�J��x։�x}����2>N�hW�p�$F���c���w�8\.��U>��M�++�>y".��B�Xy,��1���a��T�C5رs7��ꨉ.��:�΁d�Tօ�	�p��� F��lY������B4ⱨd�4r�?��e�o���K��z{��Y<N�c�p;r�{�hm�UX��`�=��\F�ע�ǎ��!����B<j�fLm��E>7�Cb��q��ޮ�.6�J����j{S�<vwt!�J�O������/jc<h��"�^bd���Oԅ�3і�:�EId��%S���C��3���F���0?�ݱ��#� ��U�uIfN<�t�Z�_���&B�E�9���2*����C����G5n�h�`T`�s�y��I�xu�R�?�/䬰0dq"$ϒv�s�#�B!#ӥ�tsgϑ)[mM��D<@X0�CCx�������wO�V�%���E����`l�x)������:�y"�4�.XTZ��V��s��Ȥl��)=ܸ��V�qډ+�y�ZćD�$�����^*�p�]���60��ett� ����=�@d�ugy��s����WzF8�P�n	>��P�BԔ�*,��)�ę�@2�8
mE*��E!�/�Yr�i%�r�JK a��)t�T6rԐIN&��"����p�[� N���0km;ww�kk�V�1�Y�����64<�
�[�h��s]�8M"8�m�&�2qmݺՕa,]�Xn����Q���аT��>6oۆs���>�q:�h��3_�@��M�3?v6���k����0e�4|��ⷿ�6�[�ǉ��0&�4����Ƿ�׏�(�d�f����N?�L�h��g���['Rۈ�ˎ��m;��#�*�ȣ��ҥtB�y��;:�������JJ뇖\t�ů䓓�;�T��EK��/y6n7����޵M�3^������As4��s�e�8�s�A_���f���ƙgw�� �m�$E�I'���5HƢ�{���"��#��I�-R3�z�Z,:b�_�'�rFi�~ǏD�_�h�͙��֢�sеob�A9˒���(��L�>C*AJ��84�N@o��{��Ȍ�e�GD�.�ua�4Vc׶-���b�Tr�A�_MWo�8!���`"�#�;��� ���"�p�죇�MɧQ�����p���|gBk�]_��W_:�q)�����YS.W��Ԫ�Ͼ����M����Uc��J���QD��84���/�z�=δDT6��9n9�મJf��%ʒ'S2�37Sm��$D�`�����@z�GI�.�Ip5A?�M����,/>��V�Wｻ�?�,���̗bV͈�ڸ+�)�K��:�g.Ƥ)s�?c+�L6��+P��ّ�ˀ�I�\�qJN�x�asC"���<���t<
����߉�D���a�����Lqv�dFEV����.)|����Qm��\'c&>�'�x<V�\�_��Q444���F�+���U�����w"St��@��vu/����+v��69�4�fs��7M�,_9�VTt|A��D�8H)'G!N����sPp��\�Y�ހ
5�3��6��IBN�L�b�
F�lFb�}l���m(/��l":�,@��Af��2�{<��ae	U)�RQ�n��Dvh�Er+�z���,PhdG���ژ#��!��6�7�wu �K�<KwۓW����#��LҬ_�}��]r�ܾc�E$-�i��?�p���B�F'-T�X�̡��C�.VL��0���*�^j�p��'a��w1�׍�@F��i    IDAT�ȏtz%j�Q�Z��$����#� _*��3
%mR�/2$nM�R�lǂ����zQAf۸��x�]��N?"+$���"�1
`¸�r'�̕מz�R�\AEEgW��Z��UzO�8Х��磱�_$^I�$�ҏ�吝�	����I1�a��T�G�	�}~����2�sU���TSU���Ýk�HӍc���������:̚5;w��������#���Csc���Wu("������,�[o��\@�o��]?��B,KXv�r|���{�ֻ����?A��'��8����s�V)��=�&�G.CSM�V�����o���r��7o�[�7�|M-00ǲcN���x����uܱ˰h��ȏkm���[�e�f�C!d)��b8گ׼����'/�j��bgΚ�o~�f���O󙫯��MmM�j�⪧�G��}����>w��T��y�ohAWwN>�t���z���g�y*
T�㨥G���W��s�>'Cb���(?簹���bڬyX�q#N=���!������u�b,9�0t�ۃ�퓤�>�O^*\C�����O�U=C<�̘��D^y����c�Aߐ�n�[~4����V���fί^S���N0T�d��ɓ�y��SiԵ�!\ׂe+O������W�LF;�?Fb<��w�R&�X��QQ��u�g���u�H�O�����]ÑU��>�7�|=���+����ɇ*�,�F�5U~�򋯺��"�p͞��[��⍴��wWW�I���7��>ڦ��<g�N:$�H�u�{��v�B9��9��%��T��Xr�|\��O���.��-x�ٗ��;����>T�C�����{��,�(�X��dL�6��#�܁���T������,�H�$$�B��N[V("��G?� �d|~w��u*\���y�U��k���Ô�tn/fN�!�^~,�r!'�<�Q+W,�E矧�i���8)����߁c��_y�?�,����Ǐ)3fa������OI:K����,o))��0� )J,�ɟ!��BA!�	a,���)1Ţ��e�.˰��@$R�ݤ�B��TB��(�_���!�%�
���4|r!8���!�vU�������u��S\ v�T�@n����=�ٔ�!d˥Q9C!B���Oң��MS����%8�.k
5rp<��׆uk04�'�y���8z��ڶu��c/^,g�={�a�&�|Ig����&����.T��[[spda�qLgy�r[TZ�M�����@16�µ��4�,���7�V��g��-�� 6ԋ��~�ҹ�i�%�����p��"��J�GAm]b���u�-�2��ۣ<�<,��ҴJE�5�����Tv��EN%�,f
RHp�J�fg�pH�� H@����q�0_Ph�PD��`H1O?��;G.]���ʫ/�w����B2��I���s����\U�Jͱ=��>��y�����A8���mum�\���}o+�{;�4�0�8I�$��a� &�NNǹ��+ͼ�*556ȃh��	����7�,TdΜ9���K0m�d�O?�{2�|9/^(���*��{�X0r�<~x��Z�T^vէ1�B��8���/`R��x�I24�; n\�1$�a�AM�<ݝعm3�i�J0Vp������w �ڧ�o`+�?�����_���]���>��}xw�j#�/d�I���[0_Fe�}��?q"�����ֆY���߽;��DC].8�Sj��Ξَ��~=��ZUN+���n�K����X> �#q�x� ���Yg�W�_K.�Ht;wl�@.�Ȉ��}�
���ˏe��ٱ��q�^�����Beтðk�f̘:	�����oH��q4�8��$Ѳy���ôY��*���E(R���g���-j���C1�B>��򣖠s���i�=>]�|��j����a����%���2y��x���ذs/�y���<$��Gu'��Ot���'�8����[����Q�د�ʶމ?y�7�v���e����I/dr�3�j��W\q�Q�	�����Pٺ��fO��3R��U �c�����ٖ�������{H'�0н=�ۑK������KJ}S�a��K��+.G[[3&�7 :��wރ��y�}
e'F	dJ���3+|�մ`ٱ���W��DpPv3؊|���� I^U.H�>���q�݉
�p����d㷒NDU�T����b$: �rd d8��Z�w�P�aJkw���I"p1�Q��9�q�I+%y�ܻ�]dT�ס҅�����ظu;�l؈�[w����1��<u��o��w�LZ{
�����B�cr��؃~%E*T؈IY��"������莝�\3�їKhm�C���[1ɤ�\F�,ɓL�AW!=f���#-*��Dao,��B����(�p#��!�j��I&J��N$�̄1�,f���x��@�4�f,Ey��5#\��Bd�0l��\",���c	$b�"�������bӦM�۱����ҥG���c�NEGT�HI����g��>��I��أ����Z|��b�2���g�G�IbE�Iu�}�,l۰ݝHǆ�K�d�w��e�(�*�#��5Zc�a,�E������o��.Ε�j���~��)L�8	]t�,҉(pT��:UU,8C�JI|]~�3YqOX��=0�X��P��|
�>j�����!0CC���Ƅ�p��k����W����!>«���r`X�=����(����_��W�b6���|���28�B��1��,U1��]4)DRf���2n�o��aEn���p���B��K麎����xU(���+�����t���
�w���>�O}��y�ir�~���C?}XM��߱s�v|�{�������o"R�����Gwc���q�����s��<��k��8�����5y]"���Tb��M����3D����K�,�*�dN�?�ށ(.��jt���]w�H2�9sg�c���������c��X�f����, &��coW'���mlB6W��y�c��#���߁�{;UБ�ńb�Γ�5!=ڇ����˔g�Y9��'��:	
�
|ꂋpߏ��W��`("C�q�B����r�m�&���$s,H'�G.��Î=��C�:Ѓ�/��\w�y/�FF0w�t�t	R�A�e�ǩ���k��9:*�GG㦉��	ګ�[&��oߊ�Q�h�B45T�?��I�V�T�d,^xM-�Ȕ�H�Buv�?�։Sp�	���x�wub��Rp�h��L+ivd�ԖZ_�ֽ�<���f����U.{���^�q�w�F�c��,�Q�s�g����e�>��On�h�ݿq��s���\���Y�ĳn�r�����X�l���c"��C>Jwy�!ڿ=��8 d���>G	���8r�B̛;��~2�����p7v��@��C<�A��|��4� �Ƶ�y�4��<���%JE��+�˘�qT@O"+Җ��V�c�-��8������i��M��*�P����L����4�P�e�nH�f�M���!�_�N���G�h>�s�>ˎ\��]����EeP:���%G.Er,�u[��gpO>�&�OW��3�#�cq�핌���c��d�oPf<�i�N���PmP.����rF]���
��~3
B�NQE���q��v�h�����x��=R�ps����xE�]��Ų�d�9��c{c?Hu�g����iw��5��I�e�GTF����L�
3�X>&��<�Gv�|-�@�*�ck��(_G1�yx_f̘�E��!��#�CC]��/��}}X�~�6ٛs��_*�>��p$&��!I����èɡ?�� *�!�d�ɘK1��O?�־�\|��aĢ���aFv�x\3�N^��V�Xy�ٹ��.�̙���w���_��906��.%0Ϙ>�]r�xGuZ��5�`����Ҧ�pQ�~
%'���j\F�ڢ<�X԰P9笳�d�BE-�Z�
ё���Tq|��c����^'/���~�����.��n���3�Bz������w��G�+?�	�Z�o�.�}�]
���\D�<��I�fD���y���/ԁ����M�3�1���G�C���<��^D�	������q9!�{����9������ ���/�ޮ}8�#���#���/��۾��߹�;������ݎ�&�ʫ>�&O��5<�ӟ��w����+�裏��^G���3�N���t\�+Dy���u͒�"A=��p4���������W�/̉��>���$��p��,�͵�2���*a��2}6�vwv�O~
s[���K1��T`M�ڮ,7���70S���S��r��FLENeu��=��h�4�}�����x��4R�"o|Sjj��Kt�/��"PSN���4<C���H����B"��7��]��ׂ�ӧJOT�*���d�1bL yP\;�v�Fl,�3���,4n��"_s�����T#96݁+�~��+Ƃ	�<3� ��������/�mw݇w�n����CϦ��o"ą<�}Q28��e_��k����)�~��ƽ3~�����9���0��,d�����ϝ~����r�+_�Be���q�����6��wUU�Lk*�R��ɮh6~:2 �����QA��Po'���HD�(�cq8�y45�#\�q�N8�(�|H���p��pw�
���FӸ)�?ɕ�H��]'�)$G�� K��r&ɒait��!he��G�i�*�x8�B�D�l*�\��2����x�4���k/�dT5�3��ř��E�d�42ԇ0SpsI\y�%h�؂�__��7���V|���^z�QX�t�6�-;;���W��m<j���ҪW1�k�/�P�c ��W��`�rE�Ǎ�#帨2��8:<��)%FR@u�Ƀ�H~9��*+5r���X.j��2�D�.�a��Ֆ2TZi��Kc���Y���1����;s��KYsI|��Xl�_�_t@Z��|M)�,D�sS��)�J���%�GQ���A�ʚ��0!�D��})ٞ1��o�S�Or���DH ���ݱ/���\v̤��W�*�:�L�?ۅ
Q��P�����p�r�H蠵���"����:�Dt�ۅ��=R��%F����s� �����W�Z�B�@/�y�YR�v��ذ=G�{ɑ2�����{�r��N:�x�ɧ�<$Nl�"��X�x|�%Ѫ>/22UY����p��#u��r�g�^t��Խ��	�g�y6FF�زi#~��_cѢ%���O��������c��W��e�^�˅۶�P�Ҭm��6oc���x���c����]'����۫e �B�������o���/~�K�&۴i+^~�E�Q�q�Y�7��5��n�]��&��8w�1zF��d�H��7���y�Y�6��O��e���x$Gc
%�D2�X����/��&*�t��N��K.�BYY6�3�$&�k���fԆÒ�ҹ��M���oU�6�oCB'�[G���
�����X�v~���F�P���ʆ���uUU�3�R�i�$iO�0]=�(r�Tx���WUL&&����nA4:"���F��N�p���"2�1�esy�X(!��XD<����n���z���O��=w���c̰'�	����� Yx]M�L7���
B�F�1���AG��y⩌�|_rO'0{�46s&*�e����B�y,��l��f�������K.ESs�{�!��H��4s�[3�N�Ķf9�y���?��E�y���n��<W~�:|����ƻ끊 \n��,T��S�'Q�*�VJ?��믹���H��_+&>��[S�������5���T����Obyz4;�>���.��������BeKG�M�`��YGD��@,�Ξ!����Ϯ��|!
9m�ȑ��(ePH'��=л��K�Q�_�1�!፥2�DP,� q��\��4�M@S�$�"��~$�4 ��A5�4�Q�b�"ӎF���P69*BPl;n����,T�`�l�Ԩ)��ix�$lVpn$�%�,V��2����z+σ�=v.C}�B�ƒQ\s�e�8�׾��iu8���׋\	%)����O|o���o܂'�yuͭ7i
�{�eDcF6��j^I#��b�UGꑈ�:9n�7���c@�D����3������� ��CIΚ���w��uC��2�Ȋ� �iC��IS�Z��d�0��BW��С�"�ڈ	W*�9zߙYL����i�,���q��k_�sYōӄ����6)��2E|�yH�`��&�0��(bC}�<�\Γ''Iܼ|�����W����|Ifo4Q�d�C9**B,D�.T���	/�?���h
�lsTH><��g���q�	�i���K�#5:$����C��'c-X��P�����}]�":4�����~o�e�g�U������ϛ+�X,>�` �7�~K7}�������!�<잙LD���ӥ_��>F�3�1I�sYt����WV�I�8}��ZQ9��#���#�a��+K���s�᷏?aT��
��|�Kp�Jx}�*��8������?/t��!ޏ7�;�~Wnǟ��u����_���zZ������=}ݸ�۰x�\x�ź&�����/�)���_�2��l����܃�׭���H�5W_�Q�	�S�&L�s�������\��q?�uj:�x�q ¹e�.�u�=شu��m�������~�7�|SF{�1h��E��	�{�m=e�cگ�Z
��ĩ�%�^��sQY]�|��x�_Y�p~?��Z��xl$���~��RMŔuzUE����r5�����#�<���w���"a��TP0kKm"�JcdM�����.�e~Ǿ���I�o����җ�w��)���!�.!���Rb^W�8i@���k���w��Y�r���[�`$�
�}��_*��G��4abk��JlV��#�� �9Q�(F�ʫ�FCK��.�� K- 8��IyE43�%��Q|�[Q���J�9�H���NŹ]���y7�n�a�a��R�$e�T>��v�:����_/X��y�g�;|���#OOO9���bgo�_;�ƚs���ӑlkU��?}��L����_���*[;���,�H�hƉ�x{�i�Y�T�< FmX�rIY�W0��d�
�b�>$G�0<ЍxlX�ٌ�vA��@y9��ŏ���K���:�����Q({Pv�1���JDD����Q�Q�y<��Hl�#;h�)�bN����ٔ�<�2"AJ5��q��f�B���\�O�u9�9|�=���!T�|��?}�Ehl�}X��;�7��P/�	_���'����������o ���S�ij�����/�oh�p5�
��r��J�4���	�DFso�H!�dzJ��!HI|(=̼�T5��JA�%7�|I2�!!alI�k�6���0.��	̘�F -TL'N����,�|���H��ި{�D�����	J�=2�r[y9� ��-"]BɈܔL�"%�����G�,CA�|��F�1D�_����H@��:���$�Q5`¹h���lȖ��rhT�yfmy�$m&gW_v�q���.:�{f#A�P�0�b�T�T� ����,��c���bÚ�@��̈́�`h�ƵK�J�Z��qu5.�2"���=���5n��3_��H�5a�:�PJĆ�%,a*w�e�HX�P>LN���
�������+0s�4!�$�0SgLW��t�7o������%,;r�TF/�������n�g?�lٲ��ȑj����?cƴ)سc�r��,Y�Y�f`��#�l��a#��N�z�i��+$�}�������5�\�c�Y������ߏ+W��cW��x�_��ߏ#/Q^�/{;��;���={�,�<+�=8:��&�,�X�����c���/�*��.8�|̜�Q�y&�-{�?a��r��������*T��6D��BA��^64��2�x?yoء�Y��q�O�	��/|{�w������T�l�HV�1�]�p�q��fdQI��k)Jx�<�L��+�BK���_a�>��/�O�H?S    IDATM�o~>��H���ӭ�Owo?���C�RE�7��y���۰y�z�/�i�e�!*�J��!��wQ1���?�H������nǁ=���5�!>�O�<P��LCE�$�Kb+Mh����g�<n<��͛���ؐ#�]�Wj+#jp�>s��#��\Dtd�PXc��V���?v.������G��6P4(�C��Q�6���w��/�j��?��r������+^�iK�p[�hR1,A�#7�6t�u�}���ʆ]�m;;Gnt>�*x�SEzGư��[:dd����(��쯭L�x2���C''gL���fL���c�s����.ˍ��]Yy����w&G7� �%C6�7HZP*��s� %Չ�!فt-t����D7/�	yET�}��`���D�rl���F�c�`��p�%K����ہ��-���8*�>�ilX���oCUeD���o7	ǟt���o�+��󯼊��̙8~���-3�͏��w ̐�~��Fe��#I��8�e?�:�,�,~nZ���b<��
v��x�� �\�t̤�#��=O�?�r�G��7G`�:��㠪�
�3(
s2L�dg���`�-���B
�m%���A��-�9��@�?ri�H���(�,$+	�~�\A�,$ױC"[	btdP(Zv�_�nT�Q��Ԫ�"!�FO�F4�#��*7���õIy���)7W��q���%^���~^�=�}K�c�)��J��%������?�{ׂ�����SjkcM5!��D�}���`)�XTR9y9+Wg�V4A�����}r��Õ&(��8�Ã����HT~"��,����CWW::�a�=��BSc���"��,ݩ���c$M;q�
���x�n���I���0m��	��(��������K.���������ͷ�����'��5����˯�	ǯ��o޸�>�v�؎cW,�%�_��h�����q�Yg��˯��{o�;��w�������~M����%D�ܲ�\�Y�_z�%<��S��>_v��6m?�G�.C*��J�4R���Ϧ��w���O>�Blʔɨp8p��G�K>�T�*Ųȥ߹�V�O��Y�0��_�"^}�5����L�=��0�hʂ����#G�|Ƶ.�3�ˢ�Ej{�T\��{�|�{�����O'B ��gu ��:��]ހA�Y��>WV����?���3��;~(�6%^+>8M��^�ڹQb�[,�T�f�TVW��B����+��8�}z~���Hr���`d@a&���ˆFE
�.����-\�X�$��n�6���'��[8���2z-�q���)�����P�ڐܡ�^�9y����{���w�!Eԅ(3��sO�Yd(�o��>դ%�CE��3��O��@e�y�w������U���̄d�˥��3���n|�X���c���{~{���ķ:�mé�h/2���҅g~c����_}����}����߳~G�����RE����&���o4��}=��X�*���0Ŋ�	��V��ޓ�eT��M�!G9�`�����9�`0�T!���,s��iSM!�
�)!��$�
�
�c�pp��;q�aU(�)���H�|
^g	5����l.��N>o6w����y�s���%�+s�g'\
3ΐ˗!WǞ���۱[j~���s1k�a��mĦ�����M��с�֭Ǆ�S0ɑx�wO"�/���H�U�]��E�/�1:�@��Yv�E��$��*�1$vYt)�yX�0��lɿ�e6���*��Ak%֪f��BEj!�0�Ft�Z�/���nJ?z���=�e�Ҡ�]���d��!�Q6[��"��4\B؊��2i��GV�,TX0��[f	߲�!�F3?�&��(̧�ߋ|:.dgF�L�6A.�9����Ա��#��(,2�ʨHgZ*����3"Rg�ň4��B����'Ld�Ft\+���z8��C�d>KzRH���a���gLBa_�̿�C�H���/�Iڐ��c$CF�KR�)�\������uD�ԭ���5>�4��Z�'��_D���f	��S^�ɐ��o|f�F��C��E�P�p�#0�?�p9ii�%�+�J��ĺ5�k��2e��?�i1O���+'ן��!���:���n���x\z�E�6�#�̅����y�ȴ�P�7n�4x��c�k>�pЍ�^|?��CB���`ƌv�ܹG��������C#CZk-m�p����׿q�m؈P0���k��,<j� �Q���[��<������hL0�߇�sg�+_��\\k��^ڀo�qf��ߐ��䢋1o�<��Ӓ�s�#N�"�,�}��&�F73�BB@�:�d���JHW���ȑ�I�,8Y�&:M~�k��#B5��JE��N��N,Y�&NRx���^|E�D�)�K��dp� /�tI�Sr80�7�K�8$�.Zt8�z1m�lۺ���E����TD�a�L��%/#B���|-t�nhj��iӤv��ljl����m���42d����>���������C�zݑ�8*�H���j�"�&����V���e%�7#P"���DY�p��������Gz,g|����e�@��<��3'5��ʏoa��ɢ�t����U.�����t}�s8ۖs��[�,���Շ��µW�xt��#�c�����]����z��yyG�:�s�o8�����%�J���C;��\5�V�bw֖d�8~�BA,j�R��ղ�)�$����Ꞹ����(���1��ɐ����Z�)I�"�/�\���o�`�V~��ɩB%y�Ud]AΞ<�io�DX�Rcq=�0s��P6��&_[]�c�ͧ;�o'���@/fΘ��;F����1��+h�6~���Sx��W���5J��݌9s����_>��LxQpQ�4^�dKL��c(�B"���
YGY��Q�1��}H��q����T���H`L��/����H%S �@�-�>�"�I��ƥZ!����؈�������,���f�X��>ǂ�\"{lHy����E�:!4���-�QA����Qr�B�~��4a!ű�yf~�5U��Y+�ؿc=R�>�
�k0i�8��D��x���uʍ��r,WD�� 6o��a�5S�VoF?.TT��}s�uȾ�a���2c2S��)��o)��2��F�s`
I��,���:
�����E)��,��$��ꈌ�l�80��yh�G�2F�4�j��n��z4�ܚ���(%�<���,�9ڐ�1��w�5
V�`$SF����?q��_P���d��B��J삷l߆;~�CI<�9C�.��b�8�X�>����[����3J6)[񿩴;v�1X�h1Ƶ��}�$x<ĒI�J�P��K/�w�?.�����u5�x�7pϏ�ց��EG��؅{�W7�ڙ5c2�2zt�������O��ضc���3f�h��ӵ����/*WnZ�A"BEo �@��>��e�3?�m[����7���S��].�3���^�\{G4����=��,|�:kB�
y>��Y9��(��(?��?.��.�ڥ��k�(��Z����Cb���D�-�C����ǟ�ގN\u�՘4�]�#׌��f�xPY��=�HDa"�J��b�+��TH�ۉ��=���S���'2f��Q����},#�b$h�ٱ�q�&���͵�Eَ�;��D��O�>�L��s�i��e��P\?B+y��R�q=ɯ��n�{;;���/ah�4ǣ��U>0\����:��1��i��Nu<����k��kTL����k��5� OHn_����L�s��IMp �������?��ӦN�H��_/M��;6v�V������Jw,�Xty��9r�����7\����(T��O�������[έ6Ԧ
n���;0�X<-��C����\���k���V|��R`�BE��!�V��E�]�Ӝ���E{.�˓;Q4U �xB��,`xh���ajL��Fo
ʦY��ޘJ%J�&��ihx@��%�hy`ه m�dѧ����T��߻m�F͈�j�0:ԏ��O=�$��V�3P5C�C�`�w�ƺ���A����F�N���_�'��9Y(�0�9��omG]�$!*$ƕb�d���2�#�kn�	9�@�P�g�!?�"�F.C�8����PU��/,�9Y�t5(�	���0>B�я
���;���
�bH�
q�YQZ�G[���(�~>G)�dʿ�+�U����)g! ���4�=�Y�#�&���(w���� �@m�[�{�h�8L"6z�R}y�����zu�>��@@�~���썣�P�QQ9�P�0�r�Z���c�CGH��a_�C9*\�,��WG���*��S������C�"�˷��j��ݬ����ƅ7�[�Q��ؠ#&�m���
��|z�h�nTW�۹�s�� �]r��֧����qy�~�TVLFSC>{�g���)�����n�~�=����زm��[��\�p.��b��OR��'��o����t����-�q<!Ԧ��Q]4,|���~�RYV,��x`���7R���}���t&�1�����n1�z��zɏ`AL�(���AOv��e�
��B	(�\N+��]5�$]~�BIfiY��'����Qz6��R:)�_[�x)��܋���
7"L������Л���4����}���h^L��	�'�� �h���#�F��!�{�>$q�QE�����%�RɌ|Q�lᠣ���LV�c8�NM!L�=J^o�l~?Ud�(br4��&��cj�O��EY�P��Q/�/�QX4��!E �1G�2�t���'��RT�����ds�԰X���^F:���E�-a�6e��`P׌�
DR�FH:W�Ǝ(�S�&�i�k�3�n��M�Hg_���Hq`�Oub�
�:�V�O}������V��!��Wm���g^�����=���l���E���������٫nZ����"�SDe;�槟{��yg�|_����F4����FI�70�� *��l8V}.�@1(aX�[����5�$[n*�w��2�G��#�4�#�%��ǲJߤ��q�:���fu �h)�Ӂ?�mi�C�\���T>�|&��o.��aCbc(�DB�v�R��ON���e.\p���[7KyA��{��{�U[]�N��W����p}������.7&N���i3��ͷ�ʕ�)z�)�Q�4���M�R���HJ^N)|�9�\h�����]�x\X<�Y��{�2~p�>�j��i����h"�,+0V�R�(mٌ��/=��*��)T�=?#'�FfF�����8*��t1�X|��0�A��`���"u�:<H��L*���ٛ�2հYQ2A�
�WW����}xo�3H�hs&4�Q��D��jk0�m<<�*�����7����Ŷ�ɇp���υޥ]L"+�0��Ûȡo�뇉YH����"�S�fn����BY�D`q��04�����H��jMm���8�S��A(�B%R�g1:D���"d�C��s�I���=�>�`����J���{ڔv�����z�T6���6���_�
^ױPR�	�,<�vu�A�9ZrE6
�VDil�>ɥ$��v�A,k������T���M�6��^�����<�,Is�:xڶs=�L���T���s����O��$66�Ұ�<<~i\	KEU���`�qG]q��+�P��H��zt
e�+�8��ȵ����G�ƓT�Q� B�Ah��=�����Z��E�:�q�Q�X%c�-D���4����d����q�]�1f��PYYcrÜ�;��>2�%��j�'�P������i=���^��GN��̜�d��a��ُE'�$��{r���<'�Y�7��8�#FZ/�EH�
�嚑����?��c~~J�/-��aQ>�ϐN�	}������%re�OC��9���g�k�j�pm-���V*�pNr��Op�p�s>W��S�^�����k>J��������f��^{SW4w�`��"jK�;�($ۛ"w^{ŧoY1�a���oZ����o\��Ưv�.qz�j���怡�Q$⦐Rl����AE�ٺu����Ns{kA�>�/�JG�0uhy�탡N�+��6�yM�~v�hN�W^�HZfk������oR�*�h|$�����ʤ�>ɏ!�"	ʡ�gn>AQ�LS2V��ys��(p�R>���K�@U��6l�C�M�d	ѱ�?χ�_|�	��hU�r"�1�|->X'�z�[���>���<�Ȕ=�j���qS�܁�hR]���*�t8;�J`�	�+���Jp1"ޑ�H�>�Gz��"Y���ǆd�pU=��ĒY�� e�2�تK��h�Ǧ�q�FM&�W� X�apq��<�r��0Rý@��/H����"\���qp������D�h��ue��cF��
�A'<�"!�2�
�p`�:��0kf\K+fL����Z�W�X�}�j`��c&���!Y�gy�[h��]3�P7�����я]�J�=�?����TP�V����޲F�o[]U��_ȣ�&"�x��K���������>U������D��W�/���^D��I�*.�b���d�♱����ٲt�f\��$�D����C,5&N�2g��L�x6��k��v�R�#*P,��e�b9xC�y�q$׽l8���j��{*�'~�$O���Ƈ�$2?G�"H^�'���$�����9Z�'�c*,��;��3��ɳ�|$��Paa����Iq��ب��8*��%��$+�.���җI��j����e8��d�速`e޸�rde'�WE*QR4Oq��B4�FR'KD��q#F�����b���}+W����&�!�Da���Z.�_������)�q����:%������w�H$1w�<̙}Ba�k��gttD�*���RI!��g���ƊDR^z�������n��ܤ�¸#�W(��~$^��m
(��-��G�d��{x�ig*��V��RZ�D>�BC���ͤ��������Ƌ��D�s?)d��>G���C|~�BR���̙#O��q��&�xg�z�z�-%�)᧡��F��DPو����ީ�w_���|ޢ���g��

��wG��'o������aҐ��;n&�����M��g�v�J���B���}/��ޗ�zbW�-����9�1�F6�$TDF�~5��[�P�B漓�>v��GEz�<��֢e5N��6[��+��q(f?�N���Q�5h7c��TT8�%7e�v6k�i�~M��j�dS�RszM��P��� R�
�ޣ
���	5������1q9���fb��"����f��F!o`E�*����"�CB�$r��Y��'ؚ���A���*J.$��P�ڎ�	ӑ�;���Ȱc�x/
BV~�kȃ����j�ʫ
ɶtZ�c��n��Q\�. �G��B0\_eRcb���X��yh̘���GB��"�������B��78x�������X��>&p'�����n�_�H}<����>��)9ʬF���2],�teC����� �t>W��N$G���S;{�L��PGR"9C�"Ǎ&&Ȓ������M)����*���-n�v�Yp��RY��C������*\�"�T�4],j�c0#�7��ņ!7���0�.D�{d��ͤuhQ����V���:g��B�Nn���3���Xt8T�s��@�Jd�"4��z'��ϰ<i**��Є��V�	���i��m 6"�S�,"U5*&��p/ ���)%���*�X�7~��Q�c�c�>�/��1��u���Bwo⩤�{��7�7�8��Dt �wq/���2���Kr�x��M�a&�k�L'00��BG��Ϙ%)1#d�2"!�>���t(��9�����M�t��kt&�M�7X�χ����cJ�c1�O�SO?˖-����"�4�M�Z>k�9� �4����7�H���؟|�w���;�p�� �H�a���6xD��d��(��
Eb@�:Q"J[�l��]��&m7��n�?C��އ��+�'x��    IDATA(�n�&S������Z�*���§�~�����w"K����d*�}O~'wP<�J&e����GBCA�G�����a��<�#FZ�]2�2Ū��};<�?�{(ɦ7ΆM�˙�ttt(����G�eŚUQ����J%�6�\R�@��ӧɁ�����6�/��U?]���&q@Բ������/_�ɳ��7\��������^���+o~�{�t�H�Q�w�ET�R�������?{��Ez�k�z�_^��ˉ�,�_7<��*���+2���2eR������M��!a2���Rc�qr�$g�CqL@c1r
d����<�Q����^	��g	�Y-���M2-���������A�$@���Q�oJwYD��aϑG9��Y͹f�%�fF���g�A��A� z��O���57Rn��6:N-��!12��%�4]�|���:dlݾ�]D��]`�X�Mf�u�L�3%ēy�$t}��E�(�Swk:{�~hd��v�Q�daP�@�N =�����\>��;X���&x#�H���O�b)*�>d5d�FA,Zyx��l%2��
?5"x�1��bc�~�z�)��:'_�¯B%T7�p�渴�f�ZF��M�b�><���` G;,T
�U�C�Gz��l�B	��'�}�$����x�V��c��m43�8c��q�H��P9������U��R!g�:->>��.���}���56a���N��X��x@�*gfU� c@�K��lt˘��Yp{T���$2�R#�ad�t�@��O�'��Le�X���'�|ȓ������E9���,�+V`��'��f����ψ�)�QA��'�Ә�9?t)�&txh5u�x�/ා=�y�-���:_+������$�E6=&��SBV�re���ݻ��O����,�A�eԉ�0�מ��L*�Y4DX�����"O=�����ફ���cW��řc{y�s�d���?8��{(�˺m���gvvf{O6m�ͦ��BB��{���"���򈢨(EB�*ԇ�H�ْl���齼^�{&	~�{������9�������}���*0[�r���zK$��]2>�{lٶE��9�!�(u��ϗ��'���Ý�Cb�縓	̵� ]�_GbՉ��H	�p8m���+�2Mk��{7n�6G�QFFV�t��E��C�
XS�n�U�^��<o��8{չ���b��w�~�C�I�=�I����7۰cnd���"��&x�7L��k��-�&�M{���Gwo�\'6�d��!���D�g蕾C#�)�-*.��s��뿆��!��⫒�KM�9���	�'^�\�x��9�u_1���Y�犽���'�y�>�,Wq��&#C��6���uK(Gi�����r⊫ע��B���ǐ�[g<:��=�$o A@��$��c��E���[{�C__}���	��}�_��}��_}p``M e�2��u�ׅ��S�4V8��?\��)���ɨP�`�-��a�/T�SO�ӆi�'���al�4_��.x�QDLQia�#qa9�}�f���C盤fɀѪ�4v�p �Y]���Y9og��S�V�Ԃ��F��c_��%�j6x���.?z�ID��&=B�����8^"���&�Sn�T�s�`�7OD��E�Z6��@ G$n��$�Q%���y��#��)P3B�,���K�?C�U$"ϏZ����i�e5M(���ގP<���A�%�x�JUbI�m��EhTo��Lf��J)"v�^�;�<�Vw9\���H�i�e�!:6(��M���>P���8�22vʻ�rEa�y�U���,�W&�b1��$@dd �e��8��LE0����Y�se���+�I�T�/ n�9
j�x�$T�es�[u0��HF("A�ߏDtLj,*�^�4	<؂�r����E�'���~|��e��i��AAoyp�#��!@S��p'˚Q�T~�v���"���K�����/X�5:�t\x	I�$Dc)e�㊯;7j5V���)�j��������WT��d(��]Y ���������f!��X��ˀ�w�"�P����<�Lq��ع]]=j=H�e�S�.B�?*�O�n���U�c�yϓ�a����s�$a�9�kh`pP6Yn.f���3����� �z�.!�J��ta�)��*.F��,𷿽.�#���%n)>'�r���@�`���#�W��.AuK�-����;�n�Ξ�!�V7�0J$�4��I����@�S�4**������>��Oa��V��L���Hd��f|�[7�������{��Y��H�Z]m��D�q&P���x2&�����FO�1i�4i:޶�6��E@���1�L����а1�a'�G��Ŕ��T��b�4.�r-/]*�ݝ�j�Cp���b�Vf�H�@V2�T����ȕ�Y�-3g����������^���֌-���
:�Fs�G�c{��8��Ȋ�INx��🮶�n��~��_!�LM���_^��!�_f�p��=����@�����J\~��RI��H�;��"cI�c���I���"���G1:��@�'�Z�Y��E����.����W8�ۏD:+���2.��C<�LvC.�K��ז�<vݥ�t��y�2����ʦ�����}�7G��#0k����d20f�(2i���{ν�/�p����Q�ʖ�}޷?�}s�`��t:[:���+=h�)�)O�74(�=�}����H`L�x��L�bT�(�S��`�f�͞�8�FDXB;3�=NZ�Xxim� 
"���O�Í�"P�8�f*.���ϓ`�*n.�Ã#���GH����D�+3C�Y4H��I}-��i��4�2-������~��KS�f�\���6a?B\Yݸ�pѡ�BA�Q+���"~N� ��W̊��i�RL�չ�h��S�XZ����<�l��{��J�&��f�Ym��>Ia�������"��@g�Fk�����F2�E,�08�</���ȭJ���"�ļ�*w�~j
$['r'X��n���L�
w�H�h��eȰ=;4��Pl�R
du6/�E�Й�e�E�Y=�\R1J�?�F��E�vc��53*]��zX�i$�cHF��#�R�6n"r2�P��	�NK+X�gQ-�m۶	���:��@��*Gِ�$S!N��|y�	V z�����S丙*�~�vf�[��|�a^<$�|R���<�%�2�/��K姈�&/���nq�QK����5�ѧ 0M:-!syC� Eb�!�N6hS��T�r�0a�F����x�7��SK��H!.cX��Tkfv�����od����3k�\����O>6�:"������8F��m�E8V�cdѶ��oL,�,��m��;x7�F~�_�����2N���f�#�M^K D��"�_[ڱ�@��gRH�_|��r���o�����J$��Hcִf4�T#�1�݁D6-y�˲���_�z�Ϙ��u�~�9�������s���"��o��$�nx{��������Ln�G]Uba��|�8�&� �P�/N�#�}КM����������=�,��lF2�fNoM�_��P�+�:#����X0����y&O���~TF"�z����Z]^���rM:�>�q�(1���l��+ϫ�o@X>։\r�ex����d���8rb�h�ˎ�b��߱pH��Ǎǔ)�%�=C#�O� �"�o�|�t���_F<��dc4Hv��ċRO��F�~a���������a�e�~�z��㡇�(���>d̅e�"Tzݘ�P/��#dZ��E����c�7���NC8e�J,;�l<��i�o��Fט�q�.�7�Bu�,�N3���X,��?a\͟/8�Wn�l�࿇_��\.�y����������/J��#9�9k�VF�|S�H�b�%��Uz�ʏ�<��5��?T��x�w�G��z�Kʖ.:%v#�-]m0����D-~�H':�)�{��Y]Q���*���ic�'-�&"�IǕ��h���T�+�54����͛B��
'V�sB�W��{yHO��E�YC�1���f�W2&��X2_:hB4��Ϲ���"���Ů��=��끧�a_ �c~�z���d�	��ÿ��m�H~7r:�&��p��6�Y� '�����␈D4(����i�����7�\���i�I�U��o��(�=7.�<�r�Í�f�"4ڋh�/'d���<��v�,�)�9"�1+���
@r�Jz����
y�Ŗ�xn�zr�G�F��"?�{&i�Z�n���ז��X*����ɰP�V�0;��:��y��)�A/;|B6���4� �,7T�a3e#@"8�x�'m����K�2���*c:�ND���h�]G$'��
PG�܅�P<:�� ���Q�� �����*P�����Rp[(����T���)���Jg>�E�L�����(�IނNѦz��Hbp�HR�߱@�)R.�m$�ɲ(��ʜ#.�~g��B��~t'�:��!`��YLz�T����D��H��Yp��ŝ�@�}�Z0n�q�|��w�7��+����� #;��JKܨ�(��Ij��.P/ş%��D
c!���`�:�o��������Ҳ1��8:�@��%�|d+T8�^XXѝp\
��H���t���e�W����{���'�V.�H&Oj�̦&��>�0�t�烳�#�����#��c7~���x������ߑ��亢�Ԧ)���������k�x�-MQWU�d<���naD$�M���hh/c10���=	�q�7���O?��������ԋ��P�b��W���
o# ���-)��{+���`.^�_��7"<�ug��q����%���Ԛ���PX@�U������Ӌ��A4L��[n��t'q�$�?2tF-�k�[�R���'�Dt��@iy�\?m��7<������º'�9�JC]��'���$I}txH�#�K�Vy�%�Y�c�n��C�����,���?�A9��w���./G�ǅb�%.�h����{�r��}t;Źx��:�`�S��S���OaO[;43��9�����O�g�a��]��T4|��e�����^Xx¬�Ϙ9���g���^�c����;w���=#e�L��d�ga�T�U\"��o��(,H�N�*���{�}�������*����[�I��S�4U,�;�h�t�x�y���%�ȋ�n�}b������y�%K1�y*��$�z��}����+0q�dX\�#��F��Nb�yh�3��H�J����������u*/�����
�(آ�������w��͟���6��Y>ů�� 5�:��p��E%�u{�	�1�	�h���"��#��_A�"�LVJ͖/;��\M\\�h�4���No�ױ��� "�� ��ѤeU�x�J��9:2$h;'�c*啯�r��0>.��q��q�2�2N������۫�dz�V����k��'�,���^\��^$�MWI,����xjT��XK�TL�	���Pp�*��Q{{�a�A|f6���#��ڌ�ƪIL�eUC.%���X��c�$-�q�'�ȡ�ŐF�ߏ�HR�ai�&M;��'̞B2`|�����C�m����&&VC~�1��eT����I��� �Mq�#�B�[��
."y��pyG���x�(V�����/�T�(��T摲m��Q��cmER�~V>7G2Z�./I�>~աݙ��<�"I;I�#
:�̗/?+N;�}����`Մ]v�Q6���J������ow�l�d YY���"���SV����C������[�Y�H�f#b��Z�Q�Eq��Z[�u���//���6��e�ຯ� W����o���}4�4(�0y�8�x�������!�y)��H� s�±$N:y).��
���{�^y-���k�Ŭ��pZ,8r�qix�	�L�6�	(�4�m�0EuW_�������zD�ITt -�;k�^�G���t�����
3�'c|MR��cC<��a5[��䉞��0i:�غ{�Fp�k��щ?�i�
̳����B�0cQ�Kp$`9J#+%`�`���c���!L�5'��7��=�Y\3�*K1i�x�ҡ[ixh ��E���2Z�]Eց�_��Ypy�k�Aa���]x�7JL=읙0��b
��Q��"@��y��"�tV��gΙ' l������;��Ӌ�������Z���h����a5Ib9�g�<�dteR�0q����;��x驰ڜ���E �}c|]�k+Q�v�ļd�����k#Y=>7�=e�(���?6mEiM=/??��o���+ ��-�J�Q��5�Wa��fR�+c� �Td@�K��wOon��y���	��i'��ň��`�%��
���ز����]��`��CC#�#�t��l���]�`J+)�Ie�ãC��|0��Í�;_�����)�Q���_��?T����[#��3[fT,���&�"�ArG��%�EZ6�Do�� ^�P]|�Ř0���a�+���G�O��h�6{6�^�
Ӛ������D-�<�s�_8�X�H!�E��I����꣹��͍q��҇�i�&�xJ�2c&��]��O=�(r���x��'��9'�/�HTH��oe/$�Ӊx&�����CF��y:�D��8�sd&��;���M��1�
�C\4� R�K�m�!�2�n��֌��	��+μþ��x�'�D�#G!���O�*��� �y�eF GAV3$C�p�@2-���+]

�s,��V*̍�[��,rt�$#��`+3�:�R��6��c!P!\bl4��dRxf��E�D*GZC݊^i�x3�U�%�U(��@R{��7�����Pbb�MH��:�UJ�����z���{�>F&�UYR"��P0 �Ȑ8(��&�q��?���NB���g6���=^ [`R���|AxK���L�|곀���Y���3~ٍEEAX*�UZVV(�r<k#�GmM�W�~�b��<�<XY ��yJE S�J⎸��r�P�H��%�q�����_܇}�����F.�FKs�MiD84*�Z"B�l�B�š�Ao�J��ȈO�~�����{RL(�4(r9�0��nB8�C_O�l8d'Mđ���������։;~x���|�r��������$i��p@�3v�u�=G]�"2<� c#/�-s�;7ߊ�~�@�E:��2fLk���jyN��|�"�U�S�.�b���b�8R0~��7�㍛��_�E�d�͟����R�rwl߅x4�SO^(�98<�l2��� ��1��q��u�l7 j��Skt���ǲ�ϖb�'�xJ�g��=�� @�ð�uc96 ����3{��(�f4L��a_��8��Sp��?�����I��S� �4��1j�b���@-A��?�x2��'/��dAǡ�s�x���k�98,^8E6"a?L:��Z�zф(�3�3	�T׊�wJ��74�M_�̳ϕ�������Ӛ��2m�rh&��G�P�����hoI��V����}��0�	6G~���J�h��C]e9�?�"6W��C��ԒY�����睄M�w"��a��x�w���� "i���y,%�#b�J�Y����4�����5KF��l2Z�=.�}��t;\���l	�GF�|��R�A��Eb�ihk�V�+��1�ѵ��pF���U��4��5p3�D��^�m��ͧ�>9���(Pټ����;��;_=;T�MY�,�ϲ)H�
Ō\�Ŷ���M���l��Uҩ�Ѓ��Ν;%��-��Qᩄj�5�\�5�]+���I1)�U����d��o=���o]�,�!J�ח�|��1�产��k����y Ty�瞶b%��j��ɧx���ʂ�)+Gm�8���)�76�����"�O�Zx�Jaq��k�~��y�1�-Rk^�ptDʛϰ��C��<�;���K��h9=�uBg�aQ�[mf9IZ�nDbYh�n@�ęg__��)ē���F�.��%�0�K/y/��#�69�	s��S�K<ud����r��*���
����VΥ�¤H���MGŜ�$�    IDAT=cҦ��7c8�B(	zye��:v��},��B��X��p9(P����.��� ��LF��t���D�`���q��ۙ3��Cl�<�3E�B63ٜ z;0��tT�����J���l�׈I�sP����d԰_�ΰ��רx���P)�����rp�R@EFIy[���DT��"G��qŐ��%:7�٢:Ok*|��З-�G���"�r[
����b)O���gVD���5�	r�Y�ιXq�r��� <�M����F47M�2���N����	��ʒ8O��Ig	jWw��I;�5��&��ֻx�U��6q�DL�2��H��R4:2܏��~����ȑO��v쀎�Kw	zGq��Bg�����+'_j�fM�*:�L2���nY���1?�;�)IJ%ӣ�Q�)Ő/��_����ɽ���;w˦Y_[�qu���	���2�Wu���\��u�Q��E�)������閭شu�����e���}=�(�p����PS���C(�8p`�6|C���A�����KE��GE�˰��'���{��^��qK�4̞5݇;��i�U6���~9d�$SKas,��g_lE����'4py��<}&���$���v����`7� *J<@4䇍z�,K`�������?Be�8LjnAw�0N=�L��}O;��}y�9+�I�����Iv���s���?���q)z���v�:�|9���_x�={&f͜!�� �׍$�PF�$��fdwI����=ІʚzaU�J�ű��o~�P8���*��h���$�Ɉ6�z)>�i^BR��k����&�,�3�/�~�=���Hq��3�Z����oy��3���nb�� JF4��	�ɐ`�c�MF��f��3٬)���|e���yweBcBFk��b���U��[��1�-+���{������wow�so|ˈ/�v��Y�g7�̪�(x�0I��`�4� 6~�8&���K/	@���]B�)+-�hu}5n���X�x1�*��,����M'�rf�,|yA&O�����|������&���랔6�>�`8�J�����^#'��֭C7�DFL��"@��g ���p;�Re��j���F���	BD�{�t�z�@�`5T-��v�i())�,(O�Led�
���J,�֭_`�7$��`�j-�?���������D��?Ƞ8%7��^y*?���?��l
V�vSB�3/ƠS�&�̊�40Y�r�+���]��¯Uo�������C]m�yq9Ͳ�,v	���M�E<ͱ���J����W�<��au��Q�ı�	��(�W3����"n�y
'�O*渇XR��,/@��'�4��3�����
�@'t� �c#����|]E�5���tP �ݽ8�ݍ��1�e�*	"'ya
@%�Η$��/��Q�@�{p���)X��Yʢ |U���3Ӧ jT�U&*J�-���hW���I7���s�Ĳ�WA�{��#�*���@W#�c 1�C"X̤�٤wf�W��Ug�;n�p�_u<��U'���#�Ǆ�#(����iZ>��F��1}�,���ҫ��ǟ��^@�x�b�li�o�_N�T����*�Ή��k̩˗�����yS�N������ ��|�A94��V�3�a����ct#�dEC�BK�����o箽�:���Ź�]��>�(�n�
�݊%��a5
h�&�2��Ă�I�b��O�䦩�⋭�a�D�W�b�S��K/��O6"�7 �V�M��뾂?��q�رe�b,_���n�b~�)l��HDp�L��Q�k�\+��=�Z�U	�ST��܃�{A�5f-\0�C�����������s��{��yx���� ����5u�`�����+W\v!���h�N���]H�"R&Ȍ�@�'������_����f�$����f�_���ضc�����,Xu)d�Q��y0�ߍuԺtGY�.��/��m���m�����R|�`{j�\ӧMŌ�(E���5��Oj_8z�Dc�:ݘ8y
>��3T�kD����@ņ���0a���8y���Uz�][*�k�?���U�ֈ>�b/�t�F��:{^|�q��<0j�y�B�Р�c��G�\Ǵr�1dd�d�d���ꨗ���B�ăJD/#;:�I�/��QγMVh�c��;��R�~ص���5�����7�� ��?���C��5-Ӛ+�LoB�� �����p���H&���<�ﾇ�˗����ӟ��֦l����KZ�8�AI.�W��\p�Ҕ��6�b�5�|��Gid��?/:��)̟>�j�Z�ݵO��7�I�'�H��]��L�>g�^��^z	��;%tgz��pFL���S)E�n�K�lΕiu���["�J��h3X�-ɘlzfǇӉŋ��غ}�c!h�
O�~=��ű�߼��9�/&�:	6*z�k1�trz;:�Hf��� �$�N�k�a�&ŐVd�(r�N�8m�L���N�v\���!\I�����"��P�	���7���c����н�3 lV׌����k0N!��ʩ��<o=�c)oQ�-��!ŚI�����l����2�J���(�q0;���W�*<���g99�����{q��~�hb$�0鵲�8g*+�E���d�J��m�%Y��o`�.7~)~<�v=Z����$�*�A]�b\˧�ʇ�����Ϥ��d��xm�H��GI�E~^�a�#M���@8�?Ō�W�L䙕�GVb;��
�剐@�V�k�8���iAɟ�GZw�Z,[r
�\q~��{�.�Q6/o�}]H�8�q�T\j �&��%�����4�}�^Lmj��Ý8�˰�Ï��/�=v��+0�i��m��hݷ�pP~C�T�c���Ӛ����݇q&C���e�<X�.�~�]r�4O����Dg�~)u�ރ.n �^o1���@v��S��ǟ"�5"-�	g�s~�qan����r�Z(f�aEϑvh�q�5�}OmF��L��m��b�6L�:C,��/�}�<��KsT˨x���Mǵk�����a��m$����Q]�F"槹�o�H�A�=�N�-Z�'7��?-So��8S4O>��Xl�Mi¼9��{�S��GסV��vʈ%����'�Å/�Ͽ�*���jX�Q��Sg�?�L�e"��U+1���h�Pǁ���>+n��YC����>�T�e�����/�#x۶�D,���O�)��� TV�
S3�e�<JJX��>t�e�u�s��.;]��>�{��&�l�&�d�&5�a��[Ff<�1/���N\$ŁdR��Ojm�]?��XB$�,:Q4.5��ªD�a��kI����=C�9�g��
`�����ká�>0��U�/������q(m���'8�12�����VYs	��>ɔw���0w� �bU	�z�|f$s:hM�d�P
���!K6�ldϤj�7������G �'�����D֎�_>�t�{�01n�J�\t�H$3��AtwFGk����'Oĺu���~a9x#��LQ�߸!{+Jp�����.�e�����i�p!�bpk�oP8}rA%�OǕˁ�$IDd�E:-����
�}����	Q[Ĵ�������*���߾	O>�<>߾z6�z<"l��G�q�8�*��@�7|"��z2�Q���l^1�Œ��̕L
k���$Z9���_�Wv�x�%��N+FP=\Yh�V$�:h�.h�N,:�L$r&t���GM��K��#�0&Ԏh�1��8�Z�w!����
�͉��wb߾v��*`���-�����@,�h��3"�$L'B�lV�8����4jKmر�]���$!m0a�T��3.�H�iNd`�:$7���,V��!˦3QX�l��!�d�.����aU��HRZj���ɍ�-�����J��dD����U"�z9u8���$�u��p�뫱������ؿw�����7H�͆
P�5��qb���w�Sze�V`Td!�\��9
B���G7���Q �u��Q�QH��
�R?��<��:�|�ұ��Q=K¬�@Z�`���ˣ�j��cɓ�
���ƾJ��G�g���Bpb6�y���_��.�?�����èÕ�_�D�O+:Z�a�����F(�E#pyq��E���;w>�l��\���� �ׯ�����0i�8t���e3���^��EY�Ϭ�H&1q�$�Y{-~��Q�)Ef*N�w��G"r�5��s&���Â��6����(i{i�6q��3���K nO9bI-λ�b<��cظy�X�/8�e�v���;wl�JL�`L^�z�	ӧϐ��]{�c挹E�8m��x��<+5�ڲÆ��)Sq�o�c�=�M?C�ǃ%'/��q����`7j�m˧��e�����S�-CEe=>�|+�V���~��hm?�G��G/�8o����:No� ��z�:��C�����Ai^x����{�&�p�JPQS��'�g?�]==�����3OG_�%Э�Į-[Ta���Yq��}���y�6����-�F��g�:����b�V�.�y�2hS!�4��	����������d�'��?�Ӄ��]����q����w���E�2}*�����.��G���*J��8��Ɖ�z��-�2��`��&��-�/��j���-Ght^��j*0:�'N�Bgu�|���%h=tz�f��!�_r*���YtC��7�52��tB�@"��;5U�b!I֦tJ��x�����=�<�Ũ�¾�	�I���l0C�$��$a�*�;HP (s1X�#2�Iˤ�o=���� *��}���v���sڜ%M��1���Tq�g"mF5{�`d��T#�X�d���⩧�a�A��y���QA���|܄|�[��I'͗E�o9��j�� �)X.��5%'��.dn(�x�����7ߒJoZt�Go�Q������1k�,\|�x��'�}�^�HX�8�Q�����*�Z��&�J�|&��F#�8��)r�"KQ8��gKSS���8(���D��|���hu��1X�[m������bZ�ō�'�@(�E�/x+�	j/�la9�(�T}K��(�lC�׊뿲V얇[;�s�����2�RCbv@ou�~��W��`ub��N�6@����Ʌ4�U4�_+�Z��|�v}���NsY5μ�Z���������B�TY��6���DdȠ*:��Q���a�ťeb#�؊a0��a��V'sbҨtJP��l�$U���K���na<������ �1?~��H�Ø�<�f�BgG+v��-3�ٳ��{����T�W��F��,��'_�a����_G?*���_*���Z|�*�3*�~�u�q���ĭǏ^
������jYT��R���絛M���ɗO*��Xm��?P޺���H&=��f�0�V�8�\u%~��;��v�v�]s�4x'a�c!&�������`>��8c%�ф�
[f���E�_�Wֿ�7�x[ޟk�^-΍C�ĩ�{��H,-���P3uj3�/\���{���a�2��������m�����=mw��̍ޞ#��:,@�v\�Q{A�ʙ+��g�� �`q�C�N=�L���uؿ����/\�"��#�h�8;�mF$2�R�yǲ�'��始-�pg�O�>��g��O?߂�>و1fT�F�'p����ηn���0>��ST�W`ْE(/)�.���ed���"(�]&'�3�13��wPZ۩�Y}ѥ2�z�'$-��9s%�u��{ݰY���>���AaH�H���}>NW1�غf�]�c���0w�Ix��a߾}(�(��3V`x�_���Y����.�iJ��r�B� ?{[[ť�2���+��K/�����^l�K��\"�>��ɓ`0���~P�>�i#X���EUM-z��D�cw��c�>���+���GV`f�D�?a6����_[���.�I�A����QQS�QH�Ğ�
��LinAEU����B"�=i�<�5)8��L����N��C�w,*���%^�c~3���arxpꊕ��#��5;�"\A�2��J,���My�d�	D� 0�>b�6Fg��vsv�eU��+V���2~��!|���F�R��K�|9�!׭O�^�P�����o�Pټ?���Go�]�Ld<N�^Ԕ��,�t�L�QVz��$�¢.8�\4����Ï?��x�}I��[��r`��q�M�Fqq��b`S���o&o���vtwu	� �G�"g:�ɱ杌EEu�Aqn,q�"���n���_�	��e"f�	<�@:��ڵ�b�Sp�O���}���b�֛�r����$@�Ͱ�̪;#�A4�D0G��?�V؊Jj=�hf�>�'��ظ*�%Iy)�7i���XX5��œ���&YR+̎R,<y9�ƒ�d��[�N���kj����lf]��� ��ڈ�X꫋q�e�b핫Hz ����s�c��/���^\*��f�Vw	ʪ�����A[{?�:4:���q�b�$Pb�`��й� {�rZث���k��
P!MI*?���e�ʦ�f�W"�������0m�!42" #�Ao6���2f��4f8=ը������bMe5�R`9�1�R�$Ɲ�,8���������� ��!�u)�~iu<a�L�F0��+�X}}=L��;(7l8�M�-�8�W�w�4*���j��'��P���F�����<�gR��_�&* �am��Ǐ����s�S�U�qS��������y�c��8�ˣ����q����ο`Q٣9S�U"�t��Y����2�߃2��_z,&w��k��������ńee��˄M���OP[� ��W��[6��"�ҹg�B�&���6D��ؽs�z��FE�r�����^FC���	,Y��],��x]8��A'� ajm�ʹ�� +����hj��^z9�Y�	��J\q�5��o~'���ǏǄ�����V������;�M�s,�B��+V���{��ދ����+��ގ7�{�;�1�K�ԉ�q��g����ab1Ll�����4��u�@�Cow�y`G$���)�>1�u�PT6E&�^u�u8�Ս'�|Z֨��R*�lV�4��"����SyU�Zu�p�X��Ȩ�W�ļ�ស�+��t'�Gq��h�S�$Ѹ��Wrf��"�K� Θ`�I��݅˯��>�<6�E5�4�TW����Ma��`o�$3&�fW���$R���+���n��Nq�>����D3�%�Y7�vh��G�y�@�tFR}�~pD�є�9*_"V���w�d�HM�׃�i�$?��8�A��0e�{��w�\K**űc�ALn���W��G��� T�n��������- �=Z8��;iΜYh�0N��<8ho���p��f�JU��s�7"�E�5�X�h1J�*,�0H�	����x�6���ح���%a��\4��f����ZV�����c΅�X����mm�����_4w]8��$�qX�9Q�NS�$��~���#�'c�,���+1���Ho��6n�(ag�
-�8�P[[�3V���� B����h�mmm�g�}�C���ql,!�
�t򰯂EZ�-[�Lʶx��������w"�Xl2��I���TN[v.��2�|��`���b��Ha ��L"Z"ۡj8��Kt4o�B�q��X�VFI�,P�B���բ��^���.Lw$���4���p!���`![�1G
FĲ&��E��=��J��c)��q�Х#r�8�����A���a��7�w8ae8���mx�g�g�!d�&��1ɊMdu�����f��r�Y3F�X��A�۫z1�)#���	m�u&9�7aɪ+17`4�l��!B�ӄD� *�Xp��0N>q6fO���?��>�B�|-����Ŧm���aG,���	�SZ�)���h�/CZcA8���hG�wyN#.����$�V�1� ����aY������ܙ-��1sCbF�M~/    IDAT���듋�e�1R_���J!B�p��|e"Tò�_f'��B��Q�q��GZ�:.Q����T
?_Y��:"FWq�o�Q *���qaU��я�qT��B����r��6��*�Z�I5K�l6�s�^�U+W�����=��RX�`�M�,����0�{U��EUV4Mk��|�@z���If����7�M���?>&j��Xp�\	 d�2It>$�|�~��`ҤI������������0�^���n������unz�$T�{d4��\�Ţ��HVWWb��f+���8�13X�0~2���o��{~�M���S&��ȉ�r�X{�z��1�18�'��dFm�8T�ԡ�`��b�4b����z��y��710<"��e��yp�٫��Ob��͒���Ic}��T����d�Tccd-8iɊ� �L�6��:�I����y�������~T�w锄6��O�0l��gV��&."v@œ�œh?܉h,�U�]�.�/~�� D�i4a4�kg`eEY~���L&6����0z��et>����3�����\�'�z�vlW�F��G3���Rj��L�e29c0���^0Q�������ޟ����O=w4`�]<�S'���B>���T\2Ø@,�:ml�֠�p��p��߅������T�H[|*���J4�UI� �,vЩ������c���#@��k ub��%Xy�X��s�c)e*%�@En'�]u.X}:\���0}�r���1o�\�u�
T�yUS��g���`��[d�e����-qa�&4���7~���}�HY��ں��[�;4

ky��j��!��g7Nx��/�7��K�������g���{#q��xRSL-J�eW�Q��X&}:^� �-zY�X{�E�3g�"��P�ۋ�!�J�QYR!�Q��y���Е%Q{��&#����qA 3�����6�%mm��5�袋0u�Y����pN��$���q���Κ���
����wJ�P<�C<�q��@�#(�AN=��*>W��aO�l�5���!?���r,�x���|#>)�b._?p��IN�Z4N�$`����]�E�ƅD�7"�+-�V4`������[@#�V�&rp�5�a�նý��Ғ!R^R��.:��;��M@0�CWO?�{����
2�,V��F�������y'-GG�0�#0[ؾ��E�A�6����s�F�|����,8��bz�c
�� �!�X�ai�f{�ғ��5����>��^F<�i+N����[�`��}D�p��08FE�$��尹+�O ќ�QN��tN��1I�ZX��2�H\@SFR+K=�<a���xz�$i��er���b牛b�Э �*��ʋU��
�l��;l
�B��y��Q1m�䁑*y ��}���_�l�T򉾅����#�.l���AuT�����ѿ�:(� N@��{�v�������?��
I5��j%���R�{�سc�X?�6+�ϝ����49qө#�[*w�sy��1��e��9]�������g���d5YE��<e
J��B�38�e�c�agx��Bd4,�ˡ�o��v;<�r��ʨ���ib��IӉ8�јd��\F�x$�9�?��@H��9ן=�D\���q�/��m[%p� �tS&����Q���#��:Y
6����ՙ�$�k�I=���w��O6b���.q�\o�-<qn�֍�6m�V��H�.�d�L�<Aj%� ��덲Gc)8��r]w��"ζw�7~��h���3�=/�����!`_��ް�5���tz�^�Z�\��9��N�d��9k6_���ZU�7m���ZT���ج�� 44 p9�e�'��G}��Eq嚵x������A�n5�~�Q����0ur6�"�Й�S�+�`(����9���{$���g_��O\�,�-*r�q\=lV��2�(#RV��pd�T�\�]tɥ������&DQ<Nkscm�K�r:D�FP�b��,��}Z�ӈc��sq�ŗ�������Ax�n�cb��ׯ�
fNo��o��֯o��.��.���J�̘,��'�m����h�1	�|�/��rm�Y��RZ�M���7~��C#B���_�����RS*�9�K����O�>���ݰ���O�?
T6,[�Ύ�������r�� 'b.ܜs>I�T2�>��,�1�ӈ�^w9fL�@( ��|�T0KJe!č�:�vO�I��Jw"��QQ(��t��iC�Pͭ|7�K�z:G}Ƣ?�����Xp�<��^d�I!�GF��E�YW۠J��he��;��?�	��oC<�ņv\�5�C "�/4~��a4��$�y""P���I�iPު����D9���%������N� 3*��	4M���.�/��"�mۢ�Қ<P)o��yK�?B JѬI6VC.�p�58�[>yq7��9U�7kz�P�g�8��x��7��юd"�ނٳ ��a��v����"p��Nb4�Bie#\�5�����қa3d��G����ڿY�i�Q�،YK�G�/�HZ5�z\F�CC>���{�������ހ�s�P�����Pk���w�yhn�Ɓ�a���Gؾ}/z��a�a�܅�
bˮ�t�֌��S��� 2z;�YZ���+b2$G?��OE���12�	�1�Tҏ���&��fۀ�q��6�l��͝�̮�n,v���*	�X����Xf
�UJ�u��� TxQ�v�90bߢ�\iK�Q9*�-> ����d��GiP�J�����+X�%�9����1=?'K>��|E�͟�gz����<�^��pڲ����K��{�삃U�Av�81eB#����b4J�:7�p ���cb���S8�N��1�UVᎻ��?>و�^���\G��K��	sf�j2 �btxP�tj��M���!j=�Y��)���m��P���0�Dۚ\B�2M���-�HA��30L'�E�*vI��L�&��p�)��_Ã?��[e��fV��S&�W-�0#�Z���CN��PL�SÑ���n��]x����^�4d��-}S-�S�����?%��5 ��:���PWUO�L�eNIRֽP�%�J��74 #��߸������s�)���ɴgl��K���lV^�lV�\*+�����#�a�+~�1c�l�v���P�Ã�J���B�*��Q��dI#�w�Ն��h�8���t�M7����=�n�"�b�?������Q���n52x��|�`�%�R�g�u���?��Ϣ��#��{��i��L4�fT���(�d���_�e?�a����"��G��!�w9�V�������������@��p�A���}��0��"f^q�*\p�%��'?E0G�������o|v�b�(jk�ع� ����>�x��P_W�M�6�W^�������Vaρ!<��32�ず;I<A ����܈D(&"����}�m�~�U�j��VS�&�g����W�_54�G��燇�_w�-��k�)}1ÿğ*M�YD��#0<��rqR!Ty���+QW[
)f�_��62H&�Ӊ<N��3	R�~�mt�0jBx��kG2BR�9!#��֫�	r&=L+C�K����Cf��k��5W����h5��DXo�c>?,V;Lf=�����ݎm;��E��JV��\y��:�JlȋC(>�}�{Qx�Ѱ��h��QIa;�.N[�}صk���hXȴ���Ɇ���IM�`�������K�n3	���,(.�Cˬ�0�K a�V�6#��3H�Ѷ{#:�l�C�i�6���Gue��+10ҏ�}�Rɷ5�a�ĩ�T �H�TZ\?�Վ����l�}����(G0�B8��Ӭ��ÎO�@_�6h5)dufT4LC���{�. ��_�-|}m���;a�eQ�c�)�q�=7���^��ٹ[�l�ҥK�h�bhݏ�Ç�?0�h�s,Ƽ�������~J�	-'b4�3G3��ٚ�ih��#�xh�C��gC
G�щ�)iY�PG�RK����q�gՄ�ظ�39���ymO�o���¸�����5F'��LD>6ϰ)�
�J*�@@r>LH M�0P���/c㼓�(�s4�O���'φ��P�r<�Rp�=*��#__>eO.4vKeC!o�'p�tr�^�d1.<�9���v�j�<�d�YNL߈��2р%	0FFDp��x pHQ �[iy�}�w�i�X��5嚣]�fG$@Mu%�&N+0/���|��MއGFIƥ���U���w�}��t��8?J].L�0�HBX�d2#T��iEiy���ٙ�SwN����p՚����R�:�M@K몪�����\Y�Hg�t���H�2�DZb�o��v|���x���D��M&8e�\}��x��?��>��	a�(�:\63,�]ND�A�[��Z��2�X�6����w��t�����V�!x�K�L����X�J֑V/��d�(^%(F�2*���b����O��:�1�N\ED�Q�\.)����X#���4�DWBw�K�}��=��>ؠ,��a��F�tz�N�x=IK����t�j,v�Ȉ�--����-c����%FG´х����-�@�I�\V,�<0˘>��_���G����-a�lbf8B$���J��av�1�P�Ѹ
��,<�)��������7�C�}�*�������SO�oh G:�1��Y$�=��L	�\}ꪰs�6���h��.Fߠ�lô�9(�Rc!�G�~�.:��W��M�,&�-�݅����/��X86Oa��i{�����{�9��e����?T6��N�/z]Rc)�x�7�:�1/ ��L�T�d.]
^�k.?�&��e4�W�@��Ц�F`f�
�NO��F�x2-v=���7T7�JtL{�h�IFX��"��'�H�6O`�E�z�y8���-)��$�J9��J*p��^���۰sO�0*�ް�dE�Vj��81���1�(�9M
����bW(���jr�q�+020$�����j0s�Q�9�#�ͼy��S���a��}Hei[4�H�Z���鈵h�� �`
��F�n�.��3"hݹ{�~�\�:m�j�xQ�)��[*������!x<�ŢI�ơ�NN�:�;�N�r:t�"���m�A������@N�%�8>���:�S�U�\�Ќ���?���S!�R��s�&��)��8�mF�mf�z�X�|��8v��&啴R�Z][`n�c#>�7��UKj┙s1n�t���z|�� R���}������L���٠�ͨ�6�6�!�}�H�|�f��М���:���R�#�^5:!��)��ҽ��<o��z�8�zfEz��1%��d@|9-�%�C����^x��l)��b5�ߛw@��`�<��Qfa� tU�u�r�#�)?����JjS�tЪ�w��j�f�aA�Rho�w�?ϼ#�L����V�y�\���{�09��H�:瞜#� �L�  �	`E��Iq%Y�,˶�eɉ����k����+{�dY)f0� �A@�<�`r�qYu�A�>������q�M������So��V=�o~�j�Z�V��}"���V�hiE2��uy"���>[?��O-��K����K�����1���c���Ӂd".f�� 7V<ę�äc�?�&BS����w�X�����H!ߕt\c�|=:13+gr<���*�)�t\�Hjߜn�X�h*���K�����?�+/��9��2��nd����fVs�B��K�¶�͉���ⷿ�5M��?p@��kd�++������t'O>�z�^՞L���D�c�mX�`.]8�5<66!�ײ/��(u�~/�pn�����x��g��Kg��D���ۧA�3�\;<��I`@PZ[_�6`�֛�q�Ժ��O~��͟�]>[@r/�;�eh���B2F=�U�|m3������D ����'����'U(��n��n�����0� j�#J��.�l�U�V��o�dm��z��o�-! ����!A�>/Cjcz-��S�[ n�㦛6J�V`l"�ݯ�U!�O��a*�Xu�����Geu���x?��bͺ���絽2	�d�H�bX�z9~��_@CM�����Z��g�ʮ��Jpx����O�;�a�*=�x�W��֎�Y�5=�9���y�]�PCn2Q�<֬Y��m��Or�ĩS��l㍛���߸�_=�S'��G
T���^|��W���%r��l��MnPt�S�I�t.d�-����U~+֯Z�yu�p��e�t7Aƺs1r�z��Q������"J��'cAnE:���)�d�ρw��/I�`Rz4�#`�E?���Akk���/��o�Q�����Ẃ��n*����c�x��i	iv�\as	�����6&JW&
�VtV%@)�G�F�MVE��)%�2�q۶mā����4�����#Gp��	��֬Y���Ͽ�N�:�^����^(ؑ-���܁�k6bx4�X��;���ؒ���S�����E �ےE9��L������\^�G�@ӱ8�s�����BB���/��1s���/���N��X e#&	6y���8qpF/C��s�b���'V��&W���±7����kE�iAyЃ`�+ ��P�l"��Q[[�ٳgk�(�����r:un��	+�~q/����7܎HڥvS$���'{�
%��0�ۅ����0��"<�o���Q	]N~~d��t�V}��h=�c��R�_6 ��k5���I4+f��Շ�4jra��R��3sۜf��Y(
d�`)�b�x.-q9�>��:⤂��6:�LF�'ۥ�
������_2b
�:���@Ne$*�]*��L@`(gEȟ��ʿ��n�L$�����`ݚU��׿�g�}�w�*P�ϔ������p�%��@�8�i�[��ce�"%���}���;���W�t����)_��V-=��Y��0����R������E�B"!�2m���������]����~�4K��:�F��5�g�q��/X�_���c��e���[�G��m]&�*�NJ�֯ӌM��R�Ê��pH3��_y/�w���p��	��BSSrONţX�h~�����Iץ��x��V�����Rd��˕g�2�N��c�hhj��������ņ�+n`���x~N2��P�����Z�7`�(�5�µE���}�]�tw+��.2Xd�)R)��g�ys-��"����υk���#X^۷�޶˗/՟Q/��e6G͘�g]�S��s���@������g?��>��O���^���$h�&҂�� 0%rG�����������3�OL��w`�����{N���ë�Ji
��3����z��JN�/���>����ڔM7ހ/}�QM���St��/����7^?����\�\k�rg'*��1o���}�'?G8�D�jQ�m��ٺi��nA��S*
6���C84Q��Oz��j�w�z��_{��	|�[��#*�{���{��C��gg%�d����#U�l�L
^KV�����Q�)`��F4՗ÒO�f�����r,�i����<��'4:��k2
��_P��>}ΈK�kȬy`�[,&�7�,�Z�y�v��o��2MQR��C���i`dl���?T�%�p޲jl���&kB�$>�5Xlj�
$G$Q���
S�R9�o��(�Mn�h��o)��v7n܀K�.�R�U3�?o16߼E���cG��a�M����d~�6�cժ���#罰 ��b��=�o?2Ӄp�c�FK}#��ؼynܸ	;_ډ��n=�^o��c�RhjkG�؊*$�R��nQ����?�#��'O����KVo�T"/��*OG�A�*=�r�Í�9�0��J;f�@�+g����{��è���XS������fEe�ϫ|%�p$��Օ��hkQ��������0�j�}�"^{�8�Ì9�0�#�ۭM �@��g����J.=dMM�~2���dˌKf�]0"M��+Ȥ��Ҋ�7oo�����    IDAT���Ө�8՚��/ʿXi��&EA�i�|�Xs�ô���k��|&L���7�1G䚐������R�٠^A�v
L�axҖ�
_�	j���f�w���<=����l#�*2Q���߯g�OHy0 ��)V�qgO��y��R���,#����v��t,*}JYy9293�q������B ����Ӵ	�2I���RNn�i�fV�|^�lעl����K:�Ym_�|��{����7��x�rRbJ����1�"Cş�V��<�yh�Ò�i�|
�i�vyuM*���
��(���i&�g�>1��Lr�%���t�����+�˵N�@�����Is��m����F�������ĕ+]8y�,�/@�k'��g۟d3c�Q�u�Q�I�J��[#.�N�����N֮]��e�>�ڙ8Ϣ��I�Z]�[�%M�(�؆�p�
,���7oV�Ŀ'g�$z�jNE�����@�Ƣ{����et|L�J�~^v�� ��y�3�=A4��tĩ[d�|�#�6�bpp@Tl	��b+� ��`l���5� ���kܹņ2ĕ�&�M�[��Ѩt2��|���<�����;�\�/����J���ݿc�����j���P����I�U(þ�)��X��,�å=a�M7ࡻoE��8��HDc����O�w��-6?��_��ڿ��?}�GT��s�wF¹GpUr�Lqg��@�UW��	8�)���u�*���hm�@Cm\�0a��{'����d�O��O>�.�cS��4}�V�%�0Pa�S��"V�i)1�5E�5�B"���Ԉ���cX�l��mRʩ`FE�4J��i1*��;-&�@�#��x�Wm�T����C�[E��Ђ���K��ƓB�S*���rܲ�f,[�C�Ja�xrYyP���'���r~n��x��I**���Y�U������X�z#&�)ēt�m�LP珽����l��*J9�x�Vܹ�.m��{�2�I�Z02J�U�u���j�9�V�N��1� �V;n�v/��
���m���C�ܥV7!
�ܝP	�v����sc���*4������ۈt*��������Å����7>��t��Ejt�ʑR8�5 �ʹ�ʺ*��0Oa͆���{�1L�h��V_5�ǧ&9�h��P�ax�*�'�QHO!�##�f��ip2�q�m�i��q;%��p�:�۷C��T(��ޗU"�����P�07��$|-.�� ŴvJSA\c��P�~����� OV��[!�gz��RTEz�.����	�;������	c�$'"X|��7aK���|����P�����pK#��=2+,�6��y��j��'���5�q��wa˖-dR9EV�?��Oɡq[��P� �W�V��s��݅��O~Jz��#�+<2��U3'��fүO�"49uݵ���ĉx�'tx�s�]X�r��E);��C{T���A�K���%�3���� �رc2��9s&��n�XLѕCY��[����uo6�X aFX��>��FL�A�T�N�^��&�!�s��xm�� ��ʟm9�[D�\)f��V|�H�B�=\;��YT���5�,��f��k�ӊ)j�2y��`��O)-��$�,A��8�K�-��Nx}D�]��������;B*1vBF6�_�9~���Df����◌
�@������f�����zծ����Á�\n�[@_�;ũM�i��gλ�9cXJ�2}�E����3�6%��|}����*=?M�fӺ�``�����蒚>��O?�ꪪp��!�?wF�����{�Sh㩳��r���M�������{g�'`q���u���tYsf�ans-f6�*�$>=�t�l$2�s��9O��?���RL��~��oz��S�38�~4wEV�0Ɵ$�1y?܊m�l鄦Mn۰~gm�ho��ݚU�jȢ֯`Eh"�W^ޭ���Ș�`�A��֊*�S��>���%�B[���w�NO��R��*�7K_�����;�pS���AD4C<�R%�7�w8y�2��Y�=U/Tb�^����UŖ6b҃�Qϼ�H�˲��}AmVl��Ba�(dΠ�b�_S�Ay�������}���b�b\eV&\zŨ�\�A�J:�@��)�m�Ut�4��)Ԗ�X_�ŋ���m�F|կ��p�m�bb,���N*k�7螿��Nd�q�5:m�I�Qi�X�@M���Bg��/[O��#XS8y�ML^=o��|�Z����X8&���p?��Av���<��*��X�o��7q��99zT�jK[�_���g�`㍛t?��$�Qe�Xri$�#
1��;��F�<�����p��4�\�1���׌A��"���Vh�O����$Rѐ�
�xБ�U�͐-?���'*fΘ����W^��E)��0jX�u��@��%�-��î�&3�\X��פW L6A?��#�3"B��+�����&z��ii�������

�{b[���MX�H�7�a��2�#;A�B&Ӻ�&�"m�4Jƅ�@y}r�������Yx=.��X�|>"�^���5���������TH|��č��*?^�Th�^L�F��N�X�^�H����9�:yQ�b�A��u0�藯���o&2�N~�:� ������x}��\2w,��1��3������X�t&Sk�Ye�w��T�q�T9q>��lX8��y"���y%?��0<L9Mɑ`�MY0l��Y�8���v8�p� �X���TX�=�y#(�}�ϫ�H��n� ��ݖ�u��1_'�	<��`��ϵ
���s���Sy߂�k��{xO�Dk@-A���:q��<�X���x4c\�ml;�o��֠��{�^�C������sʼo�a`��m6ģQ�h0�g���� �NW��i�{�Fj����[&�j�X��p�?P�Ӳh��s�n��
���rK���'^L����8��qe�fv <�ݔ�mx����4��*�0os��9�_�G��������Ú�����Ԯ���g����W�=��G
TN�O4�b��o�R�P�ؑ)Z���Rp;-�g�*��[7�h�-CǬح99:`'a)i�<�vu�'�Fgg������Ûs��3�t3�m���/:}+Xf|`�pRD�1�BN�"Q��7n�׿�uѴԜLMG�hs��D����_�w�:߉"_�"��6�w�m���U��y���@�4Aas�l�(���
�������js�deMM�6Z
�(f�G���Ȳ���栯K����l�:�N �����ÒM��$N���gކ��-A�J]=�[T�q�����׮ŕ+=�6��9�P��(]ȉcǔ��u��&2o�"Tշ"�w�����:4�ek7"PY�ɉ1�-It�y}���,�s�����k0>e6��k]�9{�����6Ta���ؾ};�;��/J0�oN�Щ�F~|��]��@���8�C�#E�����ř��8|�4�Gpeh
�Ov��i�[:O[d��φ:���&�26p�T��$��Z?�[�-��ק�Q�i1xvUܘ�u���M�w�^��7E��Z ES6nN%a���"K�MP�ŇlOH)�w	�u���bޕ6R��,��\`m6���;'x�b�uQ��K#0����<�2�,�OY��i�S��UO�м>�̃����������x��䥑N� P�y�w�Ϣ���$Eb:�������,"�)���/N����=�%'��A���������Q�la�2�r.�a�&�Ix��	"~��Р�o�{�|r�`s�u�����O�"&����:G#�D����I�}T�$cX ~��Y��i���O�8�$Hڌ���Oaۀ"_NFb�0�N��Gd�4V��kdZ��<���-f�P�K���D�a!G�m6�,�����>7�+�ˋVӚ�!S�?/��s}�����54�ɨ�����6�]���9��v��&�cE��:���{�ѣG���ؒ�g�N)�-F �%H�1y�WRK�b���Q��z%��ɜ9s��ѡ�K��O��~�@�ApZ�L��}����x��4*��deCC���:O�P�ڀ9Y}��&kH�h�A!6�$��\��m�ʚZ�v	S9��g��W�~e��P[+�Ծ�=�gr��ą�.D��j+N��,/Cmc��4F�;��D���^�NF��w�T,t������6�����wj�|�|�@%���݇�`8�{(Qp��Q�m�rF�&Ԍj~�-�Q�T��1{F��ಹ����i�p�&�#��⩧����$���@{�b4�#�4*% `�~Ѻ��+M��Z)���o/^SS�������a�[$���qq"�"��؟���8��́@Y-�vF��4���^��
x����d,�9�i������,nNsgw�\<wQ�Ҭ2�Ý�1�LZ�����A��.Ͷ�-$Hh�([ ��s�|�*��qy�ȥ`MO���7��m��5A��-[�B��#�O���IP�2�����#K���[R���vh�njbLBe��a��[V���8N\�F�p��/ES�|D#a�t_<���쇄f.Y��Ko��=�x�zO�%;�z?P_�ƍ�T%]�tQ`�c.�CVT�/��lv�t0'�;*����Ӹ��[����\�����c8G�d
o9��K��>�xN@�����b&�z16�/ ��"15&`F���G-��h㡰���݌COj�a�j��Q^*ҨًPQ/�d ���ҿ0|�X���P�Qя�}1��뇯��P�}6[�%��i4�q
4FL��0�cʫ*uhd�-�JtЄ�� �+?��V�,z9�t�2>��sӦM�.y0�g�/C=�
�@�V�>�Uf����W�cт�Ȧ2j���I+�U�V��v1����W���L&���h�������9������λd`�bǴ2�WR�VUY��i'���l��Ɖ�ްM�I;����.i �&��;�ӣϮ<���
��(S����.��)<���=����ի�u�V��jr��O^ǝU�'�g�ϙ���c^��������}�18�	3��V��g��>��t���H��h�NL^K\lڊ%Kp��m�3�~.y�V��	J��p�$c�\����W�{~555���^�{�۷+�$Oi�����2(A�Q�	C���X�R��d
�k�n����}��m�)2��@�v�ܧL+4����LҼx�� ��0�cy���l��T�V	OJ/�#�E�\�Q7S�� �a���X�r��qjtTxo	TJ������`QaX:��?��
��X�q�}d|L|j��j��2�=�M���E ���k���r�|~k��Ӄ3gOˎ���ɥb��<���$R�Z�M�p#Oi�ٲi�3�IK:r����廷o��߼���������#��w���P��x�YƬ��	Fj��iX�1��-ؼv	��4ڛ+0{F��|!;[�2�
0�ǞW_ë��a`p\	��S�@J�D�� ���l��RcPe�VG*��ZaQz���?�M[oR�)45i*μ4������*)X�����O"���
����@[����ш��fIC�kwٍ�t+&�դ�O;��m��uX�d	F�����1{.��G��]bTXA�Q�g�����\�k��U�o��D���C�l@zjW�F�鷀���B�mǣ�z~_9�|�ܞ�̘jjU�����š��]]�1��U"Z��~�������dֆ�}c8e ��8�.]���5YQ㳡��Q{k{3��E��eX�f3bb:p��{���#�t��P�Gk�L3Y�Lh��5%.���!"���y	A��"�o��V|�׾ 7�������\���	�ga����
	�pL8��e+`r�S�#�92����D���>/�98���!Jm�B#5�k6ͦ�F�?p�bxh���,�R4j+V���%���w_o�p��z�����b4*���)��PVߝU4)uj:,<ni<�kjqǶ�1�m�,����W�P�5Z�)kb'�j�:,�ߔ�� bey��#�1N��9���~��	T����q"��Q���w��A���혇+]W���֭e�?ԯ����-=�"xT���a����ſ��%ЧW��Θ���#��&,=N<&&���,�ȨH�l�DB ��t�r%��BS�=�C�bwO����ct8lsQ�����X���FL���uY0���?��L�UZ�� � M]E�j�0՘�K`�����r��}&��[��/��O>�P$�˭\N�pO"�`��	�^�%�)��y��S[)/���K��s�>*����>���Q�>o���G
���L���X9���(�L�Ο?��~��A������h�$ϖXʀa:\k�j�`�9��bv�i����W���o��R�đ#ǰk�.��c�'vR�C�߳��8�G� 
z&K��ի�h����z�o�z�v�5�9����͓� AR�,[3�*+����*�y�*�~�i�<yZA�;2�EQ9�2tϋ�0^7?'��I������������7�]�ON��"��O�g�B�Bp��UU�^�(~��M��o��s:p��	M��V��>Yk���09U�E�*d��j��OO��'�j���~ǖ���Ƿ�A�5)P968��ܞS44��D<g�)��J!K�� !�*�e��p䣘�R-�b�p�JL�*c����N8x�.v!J�Ō�b�b޸an��i��B�Lo�T��ϸ@L/�=q��2��dЏ_��p���E��V����N`b<�`����'�J8���_OY5Fä\���T���mi�����C�mz��Q�* #�$�I���PS]��{^C��~U���w&'�ؽ�5m|7޴�׮��ݯ`��K!O���aw���P^Մ��6`"C�n|�+"#��|WN�p�RpZ3�hoǚ5�Ź|��6���*����fML�С�'=]��.����7�
���D$���	�E0͢�c!Zg/B"Gc���{�Ȩ䳰��0k�2�X�#�ݣ�γ�>w��8����: J�0�-�<�3Y��>����a5�5�����ض���K.�7��1���8{��޻Ћ�����0�ZN�L���quf��T��I���ɑK*̘�A�{��q��I�r�n�dϰ�"0�{MUG6�����F8HUSo�!=ʇ�?����/�%A_����Z�|	��bf�.�C ��Y}u5�ܶ]�`߾��)�͍���4�"����=o�^�E��-�qaM�2)��x�7p��aCs�s�7�x����A�����;��� �7�Z��6����X�x)��ݏ�/���pȘrQIaf�4�i_�ڸ9��H�R���\�D۰��u�ğ|�YQ��	ndIz���y�H�
�qNd��D��y�Y���������.��!��mQς���<��Fa���>���;�>PW����GѨ��}���/jr�>)��i,�ÒmD��L�pot�TS�C��\X�z��~�=x�W�k�^1*dZ������8���F'f
9���@V�lV1$l!0�<�m�ނ��./��]���d<*�5�Y��QspJ���i7r}n�~?n��v�O?��8pR�k�fD�|-��hx	�0�A�'�B���o�5�96��y����Q�pH���S�Mf���9#P!�ɤ�x�������L50�	�%Ϡb�[�t����4��9�Y2K��z���~�c���[��rI˺�Z����8�.�d��[Q.�^�`|�������v���˗�aڴ&K��Uy�N�>1udܙD��KY��+���c|r{_ߏ�p��J%&���N��tB�P��Hg�u�(n�RѣZ*~�e݊]������ؓ�u>R�r|0Ѷs�����'?^p��y�fڇ�H:��9�����܋���cM�����7�J�fΞji.�=/�ƫ{���wQ������0$��V+����Z����]��������Ф���ć_��Wq��ۑ!]�`��Ch"���a����ER�I    IDAT�G���r��;X�ɩi�S����mؔ��"^��,F�%YlQ���97l��8�����ű��ݚ�g�G�|N;v\�q[����سw7="[~�'+99�@&�DyU3-Z��DY�n�G�@.�x�\:~ ���p�p�S�uܸ~��/\�ԃB�n�~���1�����i���ȦVL���p(���I�M�i�bي�6UP^k'��k�O����б�,^�a�yZm����`��	���\m&V�S���th�"fR'<e�F%R��04�+1mKc5\6�*뭷ށ��)�Gp�� z'��P�0Sb���)e%9��z�y�� 9=�����+�ָnUe�ݼ��qUa��٣������TK�i�#%���" R4h�0�R;�->�|_N$��ס�4J��)�0E�f��{|�q�}l�{�h«��_�����3xꩧłp��kNOGt�ҳ&C�M�H���CA5n�2�1��|�+b:��C���	X<l�,Q0ɍ�U {���J�|h���?���܆;����C�:sN�=�{N"Q̬	��pp�t j,�@�]�Uz��y��׿��������@o�,-�ɨ�sM����ă��2*4�3z���'��چ�����>ĩ��.���J�@�'cSVi�j\.�+-�m:(�y�Y\�vM���U*r��V8�=�0i��gAeD�9�����2�گ��v��5�_:�L��?&�ҡ�h�����a{���uN��-�죟F[S#���J���M�3e��s�rӅy�A�2N�万k�[���hK����|?����{M�2E�4�K��Zkd���-���LT,E�]�<[a��\~�_R��3�����kԼp�qxS4,Y~M��D�Ƃ|UU�x���MQ��o0�([�l��n���e��1�8��$���0nQ��U��/}�����D�Jl�
�90'H�}$�c���Ø>/K� �
uTV|�3��o����i�<�~6j���@:��$$1�����IgP&+���flܲYR��gNc*׺��ʪ���Q���'�rffS�H�LK����?��g�޲�ߜ��o5)P91j�����P��hc�Qc1*��͍�S���ڳ��e��Ҙ�Z�y5�K������Gc]y���^����1>��/7$Qx���a(>�M��nn�<�3ڐP�s$?��DyT�S����׾�ul�u�nB�~���J���k��?���6��� �rLǓF4g1�f�X�Z�J���?�c_��䄴��3˄�)7����Gl:.a�����Q����[o�Ï<�����)9��l�J��GM=�&Wbb:��r�|$������0v�(�� �iTW����Q��5ux��1���㍃q��9&�Mu�aGB�����/|��Cصg�M�B?��`l:���V,^��<�<��;���Κ6G����kбx-�.�Iy�ć���iT��X4o.֯_�M��	}X=�LL`"l���<5���es��ULM�a >@����6�t���p����}#���!�v`�M�l���Ѱ��%"��309܋T4��2;Bc�轤^x]M6�]�����\^O@�VάN��V�Z?�.,�\|�0���Y6�bHZpN�L;��ֵ�~H�*0Tt�5���#O�B���}��H��B^��o��8s�^��r9Ӗ�ؾ��0|؜��a��M+����طm�K��+�]�(n��U+�xbb\c�����,>{Hr$�S��-_�mw݅'RY6��`�H������'��8?55FwA�9��i8Q�,X���
|�[���o��( %�4�p9�G��'
� ����	�'���J�ﱾ�I�']���?@82% mƤ�Y'�c{��Ff�_%�A��χE���&i]^yuzzz�p���Ԅ�	�#K�=���~��	�YM��O.��9�u��c�믫�J�P2'����4��X���\2K:�)ʤ`�n�z�Shi����%p���q��X���.}>��?}w�6�s'���j�-\��w<��������`��\*��� AA�>*��D�L:'u��ɋպ�Ӌ_�e֣΃�Ny����u�X�dƀ �k��݁��*��SDsA���!�ϔz5K'�M��|�H.>b�����{����'���Iv�ړB�LW�5T�x��볬�4m�d��5統��bt��}8{����k�������_LY5��I�36�V�G���L7nڬ3����H�N�����B,6�Ѣ^Ӗ�M���gg��={�[���+>R&�h>b��h��w�}m4����ј��~Q/�(�b�L��B۷��ߙCKC9f�r�1?��s�c{^ޯ�ȴ��t�د�n6�����4Z&�PƇ� R�fJA�.<f��ñ[�A�;�����U���+@���v���zg.vID�����#4���6��l���.'8*���&7S6��0c�\$��oû�K�B���e+�N�(�b]a-^������߇ɩ���>�v�@S�\̟�=ã�Є�j��bA�Z9�9����	���qf`��>���*�W,[���ͭ�����O~���:��B�����˱l�RTV�c���p��E���@�U붠���Sq�P}��xc]�`c��!Fc��5'S��Fy����p��4<�4�+�������HCK��HG�7V�tj�S�L����q߽X�v��'���/ ��(����T���J���+K~�G6FU�[	��]紑��6b͊�rT-U�lK����O����k=�{Ty�/�F<� ��)6��{�%�}�L\7��-�PJ�E���a����b�<lN��14%��S����_�����O�B6m����v���Db
���Ŧ�n0��n�L��t�ͺ����#��.G*��_�pV�V��*�>s&ڂ�w�K+t��d���v�=���	]W{L�<#)4>��ÒW����\ @�.��0>&S��l�:\������6:,td2p��y�2W���Wl!�:e��	������aZk�L<������sKM����<�+�QY��a����_+��߄��4�O~�W4���ߋ��
���`hhP�7�8�H�`^G�_���)�n@�}�`��m���?���O
�Dyo��5k��Z%pң��)ʲ};�T�����?�Z=������6��&Rb�4-i�p���i:��+n���ݏ��O�ĩ(2�ws<�lG�ɾs�G���\�?R7�I����%����\��7�:���9t�CA=�!�ڑ	!�"1�;�Yr�x�{;%,dx-l�M1���\�M=?S�׫��ǒL_���g�3������{��;_F���~EE��x����#�L�X��NF�E%&!S?5�~<����i�f�6�}�]���lr}��b����8�𳠦7JUM��$�\�U�P�E�ǋ��h*�ة���؍F��TeЭ"�@V*����C��7?���w<��ۗ�o�[���;?����C�����ε���36�'Z�i�ƸaZ�JPT�Kඛ֠&�Pin.�A����(.p��E��Ƌ���g�����д�y�r��z1�
��	��7p>��l�3PS[%�/�򿠩�Yw��Y���3N�����}�:{I3�OPy5�Dv�G�i�b�w����4���lsљ���r��^�i5N��+��U�T���.�ݿ_��mwݩi��'O`��{��hڄ#�R6XA��\�ys��Bw/��~���;���"�׮�����au�% T�����َ̜��2�1n�~�u�U�m��X�z�X0U�����	���瑵08EE��~���I���e���p���r^�7X:�ֶ/��dT��n���>�;v�p?\�r�V/_���kĒ�GWK�i����;��a����l����N2:=��Ͼ��}�'�64����f,�7���X8n��*����#cȧ�QW���\�xN��g�a������}�h9�χ��IMs�U�^��ݱg�;'�F}SI�$P#Pk���5J�T��0Sp\CEAn1MY̢Z��;��/��<�,�P]U��<���u��?�<�I�he����}ZYĢ!��1]Z�sӦ��k�bu����8��<-vf�Ez�+W;�J�qۥ��h�o����/�RiDL)^�t96�|����h�P��eq���T��Q#7���6n�ф	�赱u>��#x��i�����'�t��NLk�Ӵ���#��F����8�|���
C��Z���@N��7*�e�pἌ��>]ѶKD��ǖ%Y@�N,���dD�k�7o��/��hluu5p�l����<uyFp��LC�B��-V�d�(��������[�38�c��ʸ�@��M�f��DXq���'�Z�LT��x�	�|����ؤ�|�]c��%;`�TgZBZ�+�*�&���Q4�������3O?+�k���R"e���"���A.�����A��L�A��<�K�]8|�]ip����096&A)�h�Ӛ��a9�R��6�]1\	3��|�*Em���?5ce�b�"aFgPYY�����V�u�@����M�[I\g��-��'>�g�ۉw�����,�"}{�2qZ �y7�H
�i���>��w��MX�h1�>tH����U�x��͵Ue)�W�ye{�Sh�.R���;�	
di `
�<y��Z>�bF�����T!�������5e�{䞻^��)9P9?�h{��C߾6�D���F��c���cC�,��spS���`aG��X�p�u4�
��,⢉�l�����#�7��qEcs�x�{͸�5�����U��QE���R�IȒG�m*�r��q;�u����o}N�S� �%bb-���1|��PIR�e��`�k4�����N�=U���ϳ5C�T�r�S,��L�U�H�bߙ�3Ĥ��F��ݨ��E!W@m]���s��K��N>6���p��(��9˰`�J���F��*���|>[�� F{��ڥ��N� ��NiV�e� \.q9mȬ$�k��f�*�^�\ ����.� ǵ��|�����p����0{�2�����iɠܙ��#ob��*c���n��@=�cYx���ŻmYt�?�+g���mO!����U�hml@]]��\'&&*y���Ī膵k�i�T���A}����}i?��Z�]�e��1I�|J���� �$\�"c}�d�h�+��@._:������]��P}��j]0l��':G��b����(EOׄPpɅ���~�b�x��R;�0׼�5m i��i��7��n��z,�>1�t��a/�_��e�>1g�9Z��9�K=�r��� ��4z�/!����{*'�x�}f���4Y�_zELAM}�|mFG��X[�tb2)�[�tM'HgS��a�=�TqF�|�۰I@��?j1xH�}b�>7\6�����i������:c�ځl��O�����O�.]�Η^4S7^��r�W-1�;��U�f��L/0}&}�����i�V���=�s�x����p0I��T�`����R� �L�`�ׯ����}�l�Y-)2^��cS�Ge9Ǹ�O���Ke~w��9㉒+`tt\���D�d6_+�mĕ�A;u�\A�
s�n�8�a�+-M�����P���;�PS�����%��)Y��ϭ����(r��jVĊ�:x��ń����B]s;��r���a��F���Nƌ�X�#b�؆��@Ue�X}�SSj]��Ob��>.�����Pm-����P����2k>��=�d#6\^��S�Q]��K)��O����#@a1�H�~���U����e��`�aq)�&O�ɨ<��8q�4ʂr���S�Y\Q��).�<2$dg��@�%E�Zg�� �̝����7������+��)��'	�L�sX�f-��[ ���脬�	��i̜� ���ۧq�ݜ��P���\WU�xxt؞���Ƚw��o||S����������Q!Pyfϡo�G?��y�Dp���eJ� ���"G:�kAs}n۲��[>ƝQ}ͼq�:<x�������?8�X,��IcuӚ,�R��᩟����d���RQ����Ռ��S��?�6�m�.�J2K���,�Y=�����wp��e$Ҵ�!gu���+Q�FP�E��,����C#5P:��a�G	V�he?-�L�Q���S����0i�)X��ʐ+��7�����F%Oz2�Y��`��U8w�ќE�>��LF�?���O]C׹#�D&�A^��/C�(�����8�I0ey����\�۷߅`����s������_``4�y�7��}2pc��R�5�8�\y�9�:/����rlزޚv�Ng��!ਯ"����oa��Y ˔ڬ*��Ͷ45����d�p��nW6�=ٯe�Ų%��f�:T5�q�?�?��_b�t�(��@�Z�P���n����:Sp[S�_�-�:�������jkźի0�߇S'9>����A�WOĵYsʂ"7��}ݍV�^Ѱ��E�>ÀӢ$�F k4L�V|�����\�z�'ى�p���KbmP4GF�d�x�d*��������怔>+f/�L.֯^�m�m�K;�Ft:�ٳ��R�e�ebM��GEy�0�}�vLG�xm�>�˲�=}��X8�����q����*ñÇ�v;0g�l�L9��ىk�Ø�&0g�Rl��v|�ￏ��a2����f�x���K�_�,~����+��S�>sA�64,��c"��v|�S�zU �4V,󡶲Ba��A6ްe>���G�C|�zz��R�>:1��gɲ�*o8p]�JV�����@JKc=��k��K/�,�T,8}��c)X��At��������|V�2C�Ã��k�9�^�M�wn�]�;w�MA$<�o�-��74���Q�h��x:����`C�^�zp-jȆ���G�!�scX1�tr`�u�׍�[�����j�r_��Ҍ��:dSq����6F��x �w̜9�sfs�&�W�:7l܈W_}��hen�����I�6�c��Wl�Q��ju{�j���#�nhdTYk�x�߱.u��;��/Y�l9�;"6Z=�("��HP���� ::�*Ś��Dh���/Z�ϛ�%d\f͘���3�$���sپ�$�5Ŏ�s�o�d�����n܈�^ލ��}�m�N�𴶦���y�J�ԛ��ԋa�&g44�������!�df��"�"�DP�g5	#41"�G���S4�tx��E��8�V+f�BW�5tc:�^$�$Yt�3�Ց?�T���O=����/\hFw��>R�rn0����w�X@����!Q����1�҄T���񕚂ߖCM�=�3f4�b!�M'Hӯ/��g?��{;��8!G>�.A��EӋ��[:����~��ǖ��3v�ˆŋ��~�����U������aO>�P>�s�� ��%4�%�_���dS� M��M�î�6N�P�`�|n�jMqs��8w��8mhii����h�&��b��Key�^�UĒ%��58< ʑU��8�-��T.w :��Oc���3�q�a˅�AO�qD��M�P��L��#_� ��`,(*�'3$-Y���atv�����Ρ�y.jZ�+C'/ �N���Å*�Y�>�#��Ḻ�k6ނ�Y��3��,A��D�ρ��N�;�6����rC�>5,�<��8�j+ي��F�a]S��[��fCk3:�.��w��W m���-�cl:�pҁt�I��y��V8��ϑ��t�\���4E��P�ŋ�R�p��1��8 i��fp�+٢�#��!�Ulq,YT�F�@EP�Lf���(֣�P�@E`�g�Z�
�'�W�����fÁ��8<^�y��q�=wcx�ox� �\UU(c��݊��_��}x��e�}��[e�E#.����!\�t�C#x�aj:�W^ݭ�����ϡ�	��~���ֶF�����him��~/����\�P    IDAT�4�r���Chi���;������n��Y3�M'P_�]�n�g~�N����06n�I�g/\�ɳ�3M������;D������U��65׉����� ��'4	�쓿@"F%�g(+��G���oP��啕���5� ����T8���T��1wv>��<��i@��/��O��Cc<�&PYU�{�ہ�^{�T�� 2q�]�3Z��҈��&�X�G�=��;N�`����k�`x2��ŉ�9��=8����#MS2Rr�5#�ƼL�/�9�;�)���ϗ�iG�σ�ݍ��r|���t5\?3Z��EW��K�G.���L&�;f*Q�ɤ���W�fP�܊5�7`���apx���E2ט|]u��N'4�EP��ieM����7������#�ҭ��u�q��e��ѐ���o���A�8�F>#�EsƎx�6�]�։񐄫|_����3�1k���߆�zM��1�S�Y�s��E���2��ҍ��~465K��W069�ǯ��T�f��(2-!8'�b�d�&�'�H"�f���UX�b%Ν���Ǯ������
�f��N�"���A_w�45�oܠk��mT�`Ww?�t^�T����6\����rv1*V�O,0��%���\ydIG����o=t�?�\�U)PQ�g������x���R���@���Z
�hD��კ�T\�̧Dm-ޜF e?OU|&��*z8�k�>��C+�>=l���LƊy M�Yr��e6%_���I1S��Bd��{��Ml�|��N�<��5_��v����a��~[@%�� �� �a_�cDmE�Bi	H�Qe�1,�K��w��1��v45��;dE���#lP�){�,��l��6o�IEgΝ֢��%Q���Ǐtօ�,\�]׆�9��|:%j�(<�Vi��zp��)L�C�q�,�	������!Lt֬y��0���i5�h��Ѭ9���U���lKR�S���H�X�#�X�es�;��px|HLO��焟����1>tщAB��=�ǣpXL���%�N��	�EҲ��Ob2�E6�W4�m�2����"o�������	)Zz���zQH�QW���� N�8,��Fr�Ra�W_o�u�@�D�}���r�����Gʘ-?�y�z5�ð��I�բ��T���^����'xP�\38��BF�"�ˌF��@%���=�J�Ĕݹ�����o���C�U����
�۩
�����z�׮��_��6fNy�O�p��y�T����ӏ~F��^���s4�@�e��Y�a�T��h���=x����x�>��.y�� N_��3��`�����~�#���K�Kf��V3[�PS�C{cf�5�jW���{�kh���N�9������u�=��B�Bϝ��}�nܰK�Ctj~�Ue	�����5�Cc�d*�NZ��8�D���p�s|lB�d藓�$1�c~^':f����*И�o`�UubaF&q���5���λ����jy�_&��y�z�^�L���N����z-N��{��������A�8sY�s.E��$��<��4�Q,��}��J��v\N�5���|b����e��rｨ��G����A��܀�����2�����cr�fˆ�W�dZ ���Zn�g/\���(:,ƪ�b��b&V�\)A2�w�*�*������c���Mmx��gp��;Z��׬8q���0K/��ؘ��ɶ��L��H�2��/1 ����6i�8�F�B@�����Z�=|�nX�N{\"CMU����*>Jm׶���p1���9t}�CVVc�x~����Yr�ݘ;kB����-�E��đ�b�z�Օ+�|�	�%˖�JW�r��F���hn����n��ތ�2;�9�}�_Q�J!-�6|�
�5�"<C���QT��a<A�~dDS��wr�nk��ҿ풹���߼����J���W�~{p4��T�P�_�+��I�Q�"��yl(�;����GKk��)T���T@39��`%�@���O�8-���r���87~c���?�ۀ�%n|>��;��mV<����}F��^�WUn>�Ҧ����%Y:���G��	.\��Q�h�L��L,6'
Թb��<|�t�Tv�_Jk�m�
q��?6Aole�P[�[��"��q���*�+�ea����|_�C���c׫��Väo�Dyx�Ոƀ��y蘵�#S����v�lُ'�����)d�!D&�01Ѓ�� ��!R1�E�߆���Zk�s'Ӕ���_]+�Zf!X� w�9�G�=�'(#sc�%9������ڏ���4�z���Wy&�6$r�t�2��x������Fl��ww��� �1�d�X(�� 5;�����G���hm��S!�'��!kg:4�3��̩���%����8j+=�v�Ξ>
���MX8w.R��z�add��`C}SV�Y#_��o�)TR�\ԡ�'kIM ����~H�퀱��Z%�Qk�#�Ԑ��(�.4�7��+�ϡ��Y��5!�d��4�'��(j+˰����}�2�z}/8@��܄�a��1�xo�߃T"�ۆ;v(���#G�Å�NE.t�����?�ɩ�ۉ�K���
����;ή�~v?e�t�2j�WT@HB�1`�	E��c��I��$N�&�%���ˍo�ǉ�8vbs?l0lzo��BeTFeF�>�����Z���͟����3M9�ϻ��>ϳ���54�	����kĲ{�N�����,��K���
���l޾C�9&�fΒ��]'�������1�d�M���\��=#۷�%gNvK��*�{���2e�4y��{�>�Zm��[G���/����J��\�a�D�18�#[^Qj�V�P=����Uk�s�dٱ{�:vD|��hm�߿�^.�\�H��c�{�>/��(�e��~õ2w�"��O=#���{��\���d��+��9'���e鲅�f�J����="��?���F�h��ܵ[~�ēr��I�LOV^��d����!�xR��A��$�9=	�*�?�" � )��@J�zEZ����ݛ��?�ȣlK#��=�K���
Y�j9�+R�e��`�<���Y��fcp�(��2�;�#��%r��s�4��{�el���.�uJ�\��E�G?�o$�h��ʖ-�ߡ ��G�}_����_�W^~����%Ke�L�AǾ��Ȩl��&�&H0�s4	�a��|�*�1s�<����P�Y�`1��0I82�/���A�1(�"�B+�2	�ς���&�D�^~M�?rLZ��e�䉲t�"�?o6ym�"�;w�����E��9��R�0PJΞ��>���O�[o�)ÒK��(ܾ�5ٸn��x�F)�E2���������1a��ʒ���2Z�ȉ3}�W�ɢ�d�\���J�|ʪ�dAN�|�ޕ�ﵵK��ۿ��{}��P�}��?��w��
�jY�O锥��K[����B
��/��P���XqP��32m�dw��h�d(����ń�>�,S��O��]�v
FŃ�/LD �`o>��	�C��ņւ�_d�1�er뭷�W~���� .���^.G�
9A؅AV��!y�����=$6=����$U�f@��	=4&vt,J�ИT ��*��!�-
7a틦�\w�uT�>�g���:m3�����ڔɓ峟�W6o�"Ͽ��DH��D��ڤR�e��E2k�"9}vX*ʕI)-h% ��U���-fT�zyHƆ�Kq�TƆ�4:D�{�+H��8c��`� -d��y�o'��q��������s�d�ai��R='{�}Sʔ�����)�6�$��$��R���p�$��
hS�d�8O,U����r��^9wR�/�}`*�?�̱"�4IS{���2c��bz1�,=�PmF�In
r��1cq���xR��h�8QMƷ���9|`7�_Z��d��ˌi��26&G�!�yڴi2{�\i��Sg��/�"��vE��w��IIuv��q��2Pm����Q$�z���E�_���Nl�I���E�L$8V*��<�`�˸��t�m�s☼�ʋ��Ôǂ9��k�d�<~��ݳGvl�̽��:2~�8ٰa��۰A�O�d� G���i�����f�o����V��ߜ�h�V�ȇ9v䰜����dά��tN�(=�/ȩs�����<{����[�[��.���ȴI�eú+dἹr�t��ܱU�{�r����[n�U�\y��>.G���=g9u�+_�7�s�>y���X(��<I���u2wV���>('�엁3�$��r�P���c��/�Kr��m[��a������cB8{��9��|�BI�gϜ��BLJ�����K��>��=�}R���g������l7,\8��K��8Vk2p�Oz{NҲ�b�q�)�u��s�c���208"#嚬\�AN���]���Tօ�2G�h����]�#��:�J|>��U(9�&�z��ʌ�]����3�n-H`�b�R"[�9OfuM��}��?�sx+׬��'O˙�~N�A�q���r�n��y�:*Є�:��B��]L�fvMg 啗x-@6�M�.�e��c�R�����H���孷�u����͔	��d�왴� k��d��y2w�|��z�U{��YY�z�L�N��۔�{�z/F�1T0���.�HT�2����fXt��!f���I��2Y~��OH�����y���H�Qv����h�x�/$�ˆ:����{����nYx�<"�#�l�-Z0����j���P)G��9q���u�"e��P-`���X���@�	Ϫr��*[�7�\8����[w������3m��;;8�����XmS�Rk�hk�5����˺����0���(�dh���>"�Ou�M7��L8��m���B�?`�^��b���-[�j�x�Y�wH �I�3}��	eB�8����ʇ@Tp���!z����-�|Z�N��g�}_�
h=T�C�<?O�G!������:t�A�Z���e�DA���12<�)�Y]3x��J��=�/F�R#� �p0ޜ�@H������k��%��z��V-�r���c@|�g�0���/~Q^���<��K��`B���.�x2��2�k�t����B'�6Z���D�5� M�@Z�G���(�*�т�8F_$a4C'��tnV
-���6A"ÑZ]I��YDRH6�y"�,F0"#�=�o�%���	����̍���u	̼�^�T�r��~}X,)KK�!۝��@�D��������:��LV7'�BA�M�$�퓤�1E��P�J5�7X
`b+�+>t�J�g�����ʗI�y9y��>�[<�p�1:���L��V!��� �O���z��	8���=��P��b@Y	���Q��\�ĨP���Đn'jԄW�5�I#MzNx0ɤ*r b@:���?ib�|���������#�H�W9��
��pÆ�Eih��ۘx�T����%�W���b�Fx�Ū����=�i�-�@�L��^��9�h-pt�t�)ٿ{�}Q1��X�FJJA ��-�[7m��<���=�+*2L���*�2���.�"A�ā?S8�&���(	�t[�m��)���o�Y�573p�j��w%��Js�	jr��i�?��::'F7ݼs�1�D�^`%� �;+�!����x2FZq�`R*� ��%Adp�����̜5���SO=���H�F��:0PYX:�dS9���C&w���شi��-H���l���;0"{c ��)b<|DB�	LS�p3�DP � ��u�86*��|�̙9K~���@���͔kG+���I�M/�:[e\[�\8G�_|`"���Xу+�Q����(���
uT��E6�0 ��@;�Nf���s��6�nzQ����tyB���];���`��"kb0�v�I���ϟ�9A� )@�j5-h����K�f�Z�<e��䩧y�B,0öT����LG>tU�����U5y|�V��~�u���Z�4s�*D��T)�=����4s ��@�p�@{P�@��zPaws9���d�;;�D�Im"	�1�s��$L=��V)�<s\�h�R��4�t��Ue��7H-T�{�A���QQ&,|�гv\_p6�Y<�����gA"�����'�y�OO��#��7�\�TV/�'�y[j#��#�`�e��"����cG�Ⱥ�k��Q��U9r���ۻ���g̡�TלLT������~X����� 6�<�Bx��9| 	!��WS�,��tt���j�z�˃ed�(����>&��g���e��b{6	�������J�D8�U���ZZ�{����(F�
�����d�R*�Y�KrvpX��Z��i�Ob�4(�r�]w2y�'|[���/�2%�7o~[��c���}�/�O�����e��QiY �+L�d�U2c�<9r쌔b�&:ȱ��qV3���(��(d=qC�z�}��n$o5"]X[�Hr�=� ���㦏�(�(��;�\��*�$o�ĕ"y�7�""U��h3�`�R�]J�+�E�l�l�V����,Q\���=HS�3b�g��P�{��`?���:!7X$c��I���R��7@+@�%�%�YupG�fui"�"AyP2�k����rh�{���du�����+VS�d���7ߔ��ú'V�D�^�Lh���h�pHBe��7N+L��		�q2~��Q�1d��Jl�p[�$&@C`���� �C�E�=�k�|��O��|W���oj"�i2Y���9�-�2ÈSx�@�������`��,w��9�G~�8�J��[�TJ��ڜ�Y3�q�N�:!�G�0XNGd�#���̮���;7�Ï>*'N���l3�TEZ��k��
\}��ˉ(�[��r3��k�_#G���շ6K,7�IT]Νꖌ����1c�o�Nm���e�ɹ@�x��3Q�7U�m[�%�#�C|�u$�A5D�̳-הg@#�
#?�"��1���60x��A�����+/��M9�
DT���1���~��ZhC�����ӄ���h4W�	�d@
�~�����'&�yL�^��^.˭����55��/�,�C%'Xo��aD
R{KS�h������G��H�!҉�g8���r�1b�!A��hN�s�� �q�u�>5�0:��k��W�we��=4$Ԝ/}�!�a�A�8~3$ΥҘ��5~(tL ���2c�e��K/r���a���L]!�2���n� �2D�?[c�/�O�p���w�b��ϝe��
:Fx�����5
s��G�pdα����l��|�]�푳}�R,�I������B�i�ul�2V������F
��H���b�G坝�I%4(��	4\G�5!��o�^0끿��=;~�Y��Z�����'_��g�O��6nܸ��˗R�5�=�0�
i�)C�<������e˨ʇ,�O�|J�yg�m@^�A�^�/}���+��[��,ी	���?��	�N]�����|���y3/\�i$ x=�=�@G�s�t�<�؏i�6x�������/�q�,Y�Hv��G��O�LΝ�:�xoZC#d��z���w���. D���� ��.�p՗R�(��"����	�ߵ�B�ｷ��?mm�r��k�8?~��ay������/�k�ߤf��FNjF[dɢ��5}�<|B��oI��&P(M�M�P@�95�C ���)(T���:����� �l8TO�C^���K�p�	�_�}����Kԯ�����d�M���v�c��=�B,�L�)��RB�����i�<(P�8	��),z�� �y�����E3%%Y�ME�[t�O��2�	�q�9&*���J&3B�2a�,�;W.�G�F&'M����}�NB� B��H�&1�K�Dٰ��:�MF�Fk��{�ȭ��ciV�� N�#R2y:�A��qɄG������(�/�'v���^�����Ӭ��e�)�hGf�1�[/�@;���u����r���H���?��
�s��"�AX�9@�#�C26:��(�h���b�xq��9r��?'������T�)�{��j=m��KOZ�j>��b��    IDAT(�νl��عK^x�U�
��D�Pu��Ł7XPޟ-�C��i=ГX�\��*
�C��3�n�&DS⟄�dj����@��^3HM�f��S��3
^?�Y�_ ]�k��-��($AA��y`-Qj5�'%&+�o�]����ǩ��EL�B�%�
)ԓ�����׀�v�F��MwR:��>B�&hX��N�?�9T+��l�0���B0�8��۩@t�|a��ڟ��������� !���N	>`��B�7�"�;�-�=��k����~�@��9�!A��N������]ـ� �<&]��K�,_B��۶1��c��_&�/��a*�(��h���G�=�y��_�n�[Pq�r��N����A��Y�4���f2j������A�9�CM/�,cE��}�����MD*T"FL�q���2DVPH|⦛�܅Aٱ{?e���}�v�W�Ŋ�]1o���ڽo���熻~��֯w�8}˔���kV,�	���L%y���Z�f���ʔ�����t0���y�19|���J���`94:(w�y�|�7�,-�����39w����Ç��A���b�C�Ԕ�BKA.�7�}s8�b��7Z��,�����k_��v��jg��s9Wn��Z���Ѵ���O����8�tͤ]��~:^"�y��h���]2c�ti���Ј�=r\��S�e�Hl9�H��z����ꕗ����d��	�0���	�����阷߼e�l۵�BY�E�/�P�Ȣ�+e��Yr��I��oj"��Щ:��z�[ �h����㠨������,^�?�6�}�t�H]�jDҔ��B�|�jiP2�F��)����Ѻ��V������N�i���$�t�D���P�8R��,�NC��&�>Īr��8���蔥��WB��d$&7����a����6{r�����kA����˺����S�P��̙3��/��`[O�z��O�}N�O��Bk�qA�tS
�Q�[k��R����$�j!����8���s���(0'j:	�3�FA��X����F������Ǐs���1���wL�!��*M'��/��h�����s�}T� /P�q
O��T2�Ǫ����Q�L.1w4e��r�g?'�wߖ��4{Ĺ�����b��Z�&�P��K\�q}X#��~�w��g�%Y�F5��%�BN@�	�%&��d�
 (<�+P�^��*�h�}��A�� t��R�2�Zȱ�r�N�%��-mU��j��\w�����r��;���S0)��7J+cO�u�ʊ	7��Ϙ=G�m��#ڇ��R�'� ��Oa�;>��gxX���L*��|斛e�ҥ�w�-�h�}$3&��>�PDt�۰�*-78��9�(-?$�.��5F���ݟ���}j/5�'�� �Z.i�	RL ����*7�r+u��?�=�`(�k0����,�ن��j�0��	����I&���� w�����(���T�B�(3)@1�D�+|fm�>�^�5� &�����Y�^�����3����-����m�-E�m�a8�]�ePLӮq��mq�,�����Y<8,����-��$,���`��<�����=g~NW�5s��L��Xl���>��u�Ql���k��1���1Ŏ�@��y��f����KD�����4n\��R�U�G��sE��Cv�}�~%��z�~�ok:�oR���'O�]�\�
O=���.ۚ�!o�Ôv%�Tag��i�B�ߩ1c�g1�[|S��w�LG�9�;D)l����_�h�첻�F��~kg�,���h	ޟX��ˉCRɉ���r��6�2ѽMo�Mǟ!s{�,A��ʎ7��f,^�Z���ɨL��[�0������.�=~3��X�_����U�����F[ܡ�{�`��uI�%��=ƹ+:zh�ԄQ%!pB<���cay�Ď_x�x@�ee<�x'י�:Wg��͈�L+5r�\�<��U�³qx6�i��Jd%U�+����/0�+4��#℁\`B�i��P
t �5m�:�pR�a[e;>1�7�
�35���R��v�юo����S�z���琾�;5��JX+�����L�]��}�C����lظn����H=Nz�����B����ro.�W�yOJS5�US�9�R��~}FEc���d	��O�jòHf*����H��{����Q&�Ŭf1g��ҕ#!�Kh<��Dl��*-�*_�]!q�V���舍�|��P�df嶊�&\��cJG3�����%�8���~�͘n���"#'C��dVY���'^�9��0�h�t��p��ۤO��U����*?��L�K��v}� 
�#���B>�������ЩT��Ca��1D�*x_�H�G������ކ���^���in�H/I�)9������^�v�LT�^4{�mC�O�K	u\�M����y� V1M���YGp����Nk�N���EP��cj�	���[�Y�d��-�6��:�d��'��Hp��C��4�~���;�������E���e�3����H���L�g�DgC������)�y��t��97����
� �_ĩ5��f�������|�!�P`���h��}1�W`qf�2�4a�m�	�LvSq�8��ǭ!�VDS&��)L�rE��T���,��ݳ�����>�����T �>L{�z��̿eړ,��"pc�RBXrɻ�hn�ҩ�=Tڝ��b������⻽給t~���:"��qqd�?)2]U�Xka�=;���E�9Ԃ��> B��iشs7����������j�X��D���&�CG�K�/����A�ìϢ���z��m����W��=�=߄e%���� ��ؓ�Ć�������.|i}=���8Y� >�u�M(W�������Zn��M�L1 �'�P�s�9���)��Ѧ�8qTF��[��پ.V!y�C����$��1(IFv�|��z.�5&oV���8���c���P��t���)��ZE}�xB=�_,�q�ud�#ڐ�)�\�__=S|Tپ��!>)Ja�Ř����2mrzԕ�;���L�"��4,"Z�#͋k���:��1+3nsQW�R��^,�+Ԫغa���Wt?����]���C^~��'�Je'�%�=�.߶?~�`�
�g�>��	��� �-�Ҽ����9�!��C�D��;P���4s�"�="r
�zϲ)Y��N��E�F����C�P�2� ��e5/6�zS����`}6�H��K��TK��l�cj��%ԧ�J�/̾H��3Q]c
zz�$�Ig�&&r�P��y�,;I@$���R�=�8�&���h���A��OT�]K���7��Y0����)L{���+���h���A�����O>��.۴Q��	��x5�� 7�7�p$M1���.!v��dqf�4f%}�lE��4ٲ�Y�I��$O@ӹ�d��hC�]����ѫӟ����5{ �Ȁ�U�]�UG��.��"�q�F�9�R�}fZ��G�|�
��U���$v���;�QQܔ�(���^�Z��cN��a�w�;�*�k6WnXXwea%��x �|Sl�Eo�j﹛ ]G�#�{ޭ�Fqr��fܚ�R�S��W�0Q�h�\�B�܉�#&��9�f���n�B��k\-�9�J=������
m�q��v��;k�#�����D���� ����d±�A��s�a��T����\��gя�&�.�@�Px]��\n'��$*	�1������^�9¡Dy��Ŕ�O��u�q���E���7M����>�ᚤugx@҉a�K�д>Z��>�� ��h��o����ZB=��Aîدf9 ZK��/��t�KP��{G���R�����|����wX��x! B�%�Ǟ��<� ]������S"��=�.��h+�;��=|��gɧ�[�p���@��y�m�JE* ��u���Vϻ �`�BxPV>��Lq� �����M�\�Ã�7"���u��+���sM�����m�~�'nct5���K��pQ�6P��ր;�N����߷���t	ȭD�\ %/���k��^P�WD*k�#l�o�.J���@�f.���ny�h�="*MgW�Z����z���*��*���I�y��"��)����Ҙ��a�~��qÿ�^����b�TF�Sy���� 6@ݶ`\e���K:���-��
�񛠕mJ�F�m���R)x�4lZ����6\�p��h\q|������v�@�f�e;Xk�~ �Y������IR�i���Ui�\�JT"���6%>��A�&�Q1�Ö�T����=��G��=�r��06���2�\�IW,�2��p4~�e�)Jì.$C�56���B�<��h_,���pZ�+¶��l�<Ԙ��>�f^���:|����O`�������`Ó����y�����d��7�?J	�2�@S�;��L����ɮcڙ@T�Ug'ŢI���o`��?�ꤋ�RȨa���:����&�bF���U�^��r,��h��F"�H��܏o*�c�|�6�^��X�(G����Q�(!K���X��Ζ��ߝL��'e{��K߃��8�hE5B���@+�;IG+�`�V|v��hV|,�m�n ����R_��Z "e���͑$��J�S����h���ap$��Ȓ�s��)8��[���,M.��6��������L��9>�0`�h.:<�-'��@���D���F*�":VR!J>�?�#���ˠW�Β^���؄zx�V�G��ߩ�k��h�´�H�:"&�詜T$(�����D������d:��iAC��"
#CF@Y��j���y\R�=�iЂ�J8V�M�3MK����0/oSI<*�а�5	���1����aW�`L���'M7�?m.�-���`�ﾭ���71>��"�'��#�B)��̸��'EY><ņ�K����s"4�[��^�y�⠅lx��F�p�Tт��t������7�!m�6�;�O��[��=�fXGE�u|,n9f
�H�1I��'_��}f�2w�-����Rg->���񑿨,�'+l Ѩ�2��M�FF��Y��uL;�(���C*�p}�|>��QyF�#{p��q�s��28�T�<���] �Nj�V�&$&3=ݳ��T=�:��q���g�Ƞ>�&b;?�r5��̫�����l����Z�2��[����yS3'��^���1���k�k�e��?ȩ����rV/KE2	��Φ&e1���6sY���~(���a3o�v��,�=�ϳPy��
����}�^�����ٗ�tLI��p0�+��`9|�&w��>�i���O�x�٬� �I����p��g��XәĤ���ۙ۟W�:3����/
��ͧ����׶7'����D(����i���RʈB�a���/�^+n�Z�Hyh	J��ס�4�������n��X�b�P޿mZ/�8���h�2��І[�:R*50��S���C�$'-�$���HV��8���0�4�#|��q)~�e�Kq�BwM+˭�r%���Z�-���������?bW���C	S�o>	�\���-mp�S�����`�p��S"z���3�e��@����b�B�ʀT���@���I��q@��7a-�E�3��z��s�nq_v7-� ���uI��"���W�P@R1��e�b�@HG���]{�10XD�U\�~ *�uL��wB�"p��J�I�����Y�M]Ĵw�����{�����@	 $jP.ҭ�
��]z��������5dӜ���j&s�$����j���lu�����Ź%��t�koow��x�X�H�Q��A!9�	��9~;v����;�D�0��'�8݀,kGZϞ~2j�Y����mߞr7��NPr�=�;i7~&����mD~ZM�)���X�� M�i�:T�Vp��BcA
\qrr��#q����q]׮��Z�O��KTS산��e60�&јx���L���O�sXj�/�Nv�/-���T%�D}2��3Kj^�N35�xG֪�/�)¦��M~�&f%��s˓~	,���)3���ȉŐ��F�c-�U�C"Sb2�<���N�Z�"T�s�O�_�G�r��lw$05Bj�s�Y�������l��}R���7&��Z�����Muᓃ�/��'���<a�=o�����w�rƁ׍?o�G�S�3#�3�&Ӑ�����{�\�� ̴d}�BH�����t���)xq�,�x���9�����6��"�P�����q'�i�R�t��)!�Fi,\��\1M�^bq�P���᭖v�����,�{��Q��n�A%9|���0��W��B�Cز ��U%���en�QY�Vê�D��*��E(�*����9w���M��=�`�ƒ��NA�L��cP�?!���f���Sϼ�8��R����Eq�F5�� F�t́|!,"�rCa����?���ږ���k鄦T�uV֚=�$E�7�|\S��m�Z�� �e���QHW�k�"<�Ƚ��|Ւ�W�܃(�aǂ��p��]-��j�.�}]@�"(�COgl����uK�I~�裭Xz�hjd�'�b�����fr;��۾l�y\��>�L0|�Fٕn�k�m�ws��o|``H�2��I�w��j���竆�!����<Λ���$����xL�8�kʴ� ��$D�;��N������߹��R����x%Fb�Ǿj�o�p��)��?���z��_O�LÌ���K�#��3�.8�͘*�����MF&Op않;�T)�j��	#�,�iSR.EJV¶�O
Vq+�6ӬkF�?^�gG���tFsГ��VG!�S�;�Q�Ш�4o�����[�����3�ʂ��p�
�@㞕L��dh���n��/��c�w,#��NP����xW2�R��)(Y��9�~����EθPoO� ���L~U�|�F7�9�&p���YR	��ؐ��Sbs�-�Z�c���.E.�g�,̤=�g����	z� n ��c絣f�xG#!?eˡ��g�mp?��J�j�D)�C���[$�:���!�!��6ƪ�܌0�9iL��&�k���U��0��"�a�b���ff|���	�(`��?r���_�Y
�%�h�Q< db�1&��ܪ��b�<���媲;H��ca�<iR��I$���)2�r�y`!a=	������3G_!ޓ��j�'���ވ�n��놂���Q�c��ˠ����G\ N��J+�����T�[	�d�Pv�����/�B��O�E��I������WK*���S�L�f�1{�*Y�}9;���*���f�����	�~\$�ߩp��ۨ�������ď�����zR1�u�������[)�v�ξ��ΐW�������X�J�
n�����&*�^�]*�ݗ@<�v���[en�
�u���S4;ѻH�,���O�,g.W?C�6Va;2;�T��o~�ك�Ӭ�MH��۫gJ�19�p(2��L6Gz�A��I�rB3�|41�� �B\O�y��E�R�xT]�~i�+�ĺ�St��wAUw���� ���Oj�I[G����ݮkT%J�	 �S9b��Qc2���FD�Ӥ�1l�ٔ�h�+�z�5ia��Q2��)��zj��
��?Isp���i�#�=+H��!���}�A�t�'-�0D���[������e����}� ��3�~H0�i��06�_Nr��H��o�_r��E �+�T����oϴα���E��Ut�� �q5�f�$i�g����I&�磣iB����]sż��9K�.��IFbb�6H?���1P=H���i�<I>���)å�y�إITlqְ�I���~.V�j��|�幑	����8��j�0�㦡�?��C:ԣ7����rH5%v0Q�J���%�T*�+�,b�Ij�,��U3�x�\��m�a\��|�de���t�0��VFz�;ۯ��X��hsӮDQ���;�	�U�eA�՛e�ؖT��X^ֲ-��|����q7P��ʀ]�ʗ\7�"�J�����4��v���<نt)������*tv�C
�FD���p�����@?SY��#��a�M�	52�����Huġ���Wi�u��*��Z̃��C���pAr#���aH(�8���Fwe�i���Qi��� l�AN)�U��W:��>��W�c�ߎwg��	T�M�N��U&J�Tz���Y@�	�x�_�/�"��LU�9��FF��@�	��５T���˂~[�*��_�0DR���}���MV�ϊ����������b���R5�U��A狰����	�w�H���݇W�F<��cb���^*�=T���O�fƝ�+q�C�/r+�Z�D�
�"z�<خ����DT����pV�a�KD��fb�/����u]pV~DE�n_	~���^4|"20�m���)�>�i�)���̅!ު�X�J��A��Fn�L�]V>���U#��D��0Y�?� }7/߻�oE5��lg��+g`��c����ކ������~}����C�u�v�XO6'ڏ��]؁qy�����$\07�9�'{.�����k� 9Hu���2�9.:�fs1X��+;�� ���WחP�۶i��_�,�@f�<���)�:(�f�EB�o��]�p����J7׽���w�ڻ�w�(\3MV6�41������d�e%����M���F�ک�$��~o)�W��W��L�����/^�oN�g����,�ہ*�mR�y��c(t�f��K�!��i����D6�9]Kr!|�Ud�4�!װK�,A���8QQy@.����̠R�}�⛔���Zq;�&K:��8Uݴ��\��wĀ{�N�d~Y�j?Ia-)��:���52:
4��O�?�b`Ȑ���#��x\��n���)^$��2�I;�79<;5�u�Y>��0�w>�}Y����HAt�L�QX�Q`A����v�Mlcf�'H�ڕ����%�0��-�$��5|=]��G��@hw
_4e��Ip��ΰWy�fx�d?w��͌�A�Z��I�Lv��D�<����ט�v�\)��/S�0-�Ԟ��~)�l�#Ӡ�#Y���_g�¸�>cF����k�ym���h��:7�,tM���>*H�_Ⱥ�qm�u�}�=ά�aP.6h+�;�r�	w��j08���@��U� �L8Vx������P��8�M��$kW����F���j2�n%O�mN��Z�X�V���y$H���3�!'�J֪��F�
@�ϱH=�Ǧ�8[�՝�Yhw1q�Ϣ�תg���i�ىg�y ��;S@c]uEk\<�	���Y����b��q�l�0pZ���u�!Yܹ��gO7K��z���J-?�!���7��ʚP �T峰}�l�Y���<�^�������o�����!-��_����J�K�fu��H�iSeM�66����߲���F-�U�ϧ��{Ψ�||�M���s#���5gg����Bl���n��e[�C��}�xƷj���T�@JT=�T'fm��jg�E�o�u��nVV��S0pމ�32�3ՆSW[,�(���G4�5�����Z-�'��5ԠEv�Fj����{��z�F$�~���o0x7A��f��$�5�BX���b?��3=��?�����´�;�:�O����P��9d	u�::cE�ٗ�Q�R��X��UXsG~���-9|>��1��W%R�=�����[1I��C�Q��n��Cb��,Z6��e��ZO���+����7ئ��p�߉P�I���La�W��G�QO���ROO�f�$2���$)��9?�Y$�1���o�`'�i]Z�`�����}�\o;/��-�%]���@�
���T���	i���oz�R"��g�
��?x�tz�D�u��f��}��[]241PI�'��������k�����T�#�,w4U���o��#��BIz��X}Q��԰��v��C�M��XD��i}�C�ՎDf�
c�	����JN� �����P.�\��ݾ%kv,�4�@���%�� cU���Qt�tސ�/A�C�pE�^4%ޟ�A4nT�`�GM����L9��L#�:��������@��Lk]��� �"�⊿A
J�F�9��֬H8��lRݲ��r
�W�CX��FA��FDR�QVG��Y�#3
P�H6d����W ��(-��N]ϣmV��ך��&�p��ء��m
�u��hp�(W�E�lo0��믶�(�Z��	�<��+̤�mMä����sQyPR����~&�H����V�o���a[m���C�́P3�5�f�l@�@v����	Z���\��:Q�cl$����=<��b�x,6��������3����� r��k�_"��V�T��6?K���LȈŝh�G0w0�%����1�lM��'խQ����IQA�G��_y�׮z]�|H��v��N�[{@h�3W	���jLP}�%e(?%Al��P���t�Z3��Q���
ϏN�B([붬���p��ⴉ�#��Ȱ��tXf#x���v���x-�qG�{|�d���zv�����&3�!�	�n�?c&�ns'�bgt�R�-W'ZfYX�<c7�����MB��:�3�{R>eebb�	��7��ao��00��c��p�p![�EoR�-�7��"�#�pq�%�#��K�pr>'$F9�w�XD1� ��[t���bn��s͝�|gٲ��U����WR��������4�g�	h1u�E�L�P<Rl���bm�R�9"��d�����Ԯ}v��u����ɔ�Bf�D��t�������@a�Ϭ3}�կ#`!����t�����k��k�X�:&C��Бf���	m�sV��4+��A�Ҩ�\	{��Wp�����k�^�QWXl>��)/kN��NH�wd�N��P���c��SFFax�o|h� � #Sz7���x��Z�ķ�
uN^��<:�:=�m%e*3�*�O�J�׳�yG V���N����PÂ�̉!���I;1z����c�޸�E�����p�!���~���~�<�FJ#Fd`pp�q�"���CGr����Z���g @��F�"�-&��:��2�-m����ӂ�ip�Uj2��*F;�����k�H[ț;��4�{�Q�*̫�_�G�뀒�̕ �.3��C̓�,�n��I6����$�� 3��D�~�N�I����t�i\�DE@@�ss7��FDؒ�P��	�i�ڰ"<�#��Pw�sW�������#B����L����O"e�M7/��d��2�z �&}m�{@I���;3��([�D1��;�XӒ�v"�L�ƣ��������l�OK0v�\�������nX	���UR/�B�`��sCO|������-_}3�H���a�*-1��|�
��T�Y Q�C.@|�B�~�6'�27
��<���C��~H!$�i��VB"s��83��	�݁7u!A���ӗҫٔ~du��)l��d��"	��.h���&}���w���}uOu��{�����Z�{��O��M.§r;CTr��C��W����ϓs�rz� �|B�q���D���B 펵��̃�i�L�༷�� �v��L���撸[��ի���`R���[|ӽ����WFղ]M��f�G	�BB��m�c�D�)f���X��fG��YY��,vhvtZ�4/�o��	ٜg]���)�,~�bU������9�u���@�#�����j�އמ"�ҫ��O��}ݝ�����ZWt/'�b�4Ⱥ6����,^b�i}�!�_iI-.���SV���#���w�n��i�ӊqī`���p'��n�,4%ۆ���`T�@vV�]T|��k ���sؐ%��|�u���M^$�ة��C�)�ߊ㜌^��n�ɴ׬s�zx�@޵�jM�o���i`׶M��E�� ��nmNԩ���e��FVXӤs�M~��T�5���4��ʋ�������oYY�\�n�>����W___M�~Y���u�J�����o�@v���`KᬙR�~?Y�MKʦ����B����t>j"��qGM��{���m�R�y��rD❃@jX�7&�G>fj?I�� ��NI��F��s]Z'b��\w�ٜ�mS{ݙ6l�(�
;&��Q�7.�>��=�yP�7P��m�����׷�Z�����=\O�)�Q��ʤ�zsMK��$s��@�$G6<'N�VB�Ce��uWS�5�����-��I�Z��~��F��B
�)�;�#K>��%{��nQ{y���	��
'���BC+�X&ƞ+[�/�����:��|s��$Q��m�	��(�E�2v1r{m�,n2�[g|�RK�w��t�K<;	�r�Л������I{�O��e�����[1c��s��E�F��M���KU�*��k��!7�0/���*�d�[��i}<�0��κA���L�Ǵ��!�/hw���	kJ��	��ټ'#�BM�t=��m�(M�y&%o4�r�/F�@-�#�W���7�P�I��Y��d�pd�@{Q�EQX�N	�o�4J�La�)SW�⤀n�r��`tk�1!F���8��<�V�IQ)�{��o$�6��v��)i��)!�k&�S?����s����@~ӆڞ�ғ��_Eȓ_�,Ū��L��`��2���a�_�����!�3^Rb��R���+�^3��4(�N�l�(b�m^���Z�X�/Yf�R���ZMNX��R1Ά!H���U�n%VFBP�׷�D:U�������T
��聃6Θ���OYZI3v�<ֿ�g�)��K4;��IX��0�%��΁�t�R�;ق.�[*�1l@�<.p_qG;HI9�S@0�T+�<���Ì3��������(�-���gp��l�|@�`VFGND�6��n|���IX�an73};�ij%pbr��ue�o�՚5=�.[��7\�uh�E�9�,��naL�5T"�7n�&������̊�yL�~Ŋ��w�|���ȎW�W�t��? ׅ�a�x_����!m��������\��gͣU�<�4�0cD�����t�Z]/�̮Akʼ���|����^q�]�_A+A\�q�cc��+i���Vl�B�W�\�~(�0yy���~q�[���aZ������)��=�D���6�����ҫ����O놐q��1�k6J�k=hnu�˽�/q*�E]q���K
օ����&�g QOo~�>��A��&���NO���o�����;2=��2~��$?��[�/���������<��S��?��J�l���O?|��wM��q0��3q\�L��k�s/�8o�oJL�U���%1�������bE�x���[��������������A�}3��B�ǿ*D_u�s���a��g�?�)���Ӕ��e�-��PK   ���XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ���X����G	  ~.     jsons/user_defined.json�Zko�8�+���)����|s��4ؾ���.ŀ���XGJe�EQ��4=�	0�E�ɖ��K�s��y��*Ώ��M���b�*b6_̿�j�*��'<te�M�[7�����_6Ͼ8f�gg��u�7e�
��Xlʊ����=6?-�����b7���XG�_o�b���s��s�	�2,�0�3dAox�1��r7�Z]�{Co��]��R����	LC���f�)���\�1�*>�sW�������y��<Ym����q��4&��(4�n�������� �a�2�b�yK��y]������ܬC_��t�HL@'R���-�Ͳ�ʊ��Ֆe����q|<���F-t۠sm��z�o�ߝ��ы/[���z��G�f���7����|7��P�������Ǉ�6�����UE���.U�U��յ�^��f?:��ޅ/�����z��:��	�t��dr}�]�ʯo��������#_�6�t^����n��6����܇z[����W������	ƦY�����F�s��T���3�Q�,�*����|4NYĢ���AH��c|Y��|[������Oq���5��x���[�f[�i@���y̘S�3������`E̳< O�j w�+�� Dΐ��Y�q���4x/Uhk�(�7����|V�L��.d�9��ec�ݿ�Ĵ�,P��b��d�L�Hߤ�C�ܽi�a�)rǱ�B�D[�y�B�-`�ߥ�e��7N�Hr!�Z.3�W�U=;-�m����U���G�
�a��,��E�!s�H�=C�U�]����7H�j�����r��Eb��,%�f��A��2e6�bhJ(��5G�Y�2�8��p̪�0cH��V��z���A��9�/�Ѷ(GB�t��rR)��_>�߿~����-��Oߜ=����M�7�,nb}H�֓`!��^Tl��I��S�1�$�]��۠�/����@/�Z�m��I�Kދ�ژ=x�9�ڴ���)�Aۤ�Ӽ	��mJ�i���~�6��4�_�~�6�\���Q�������aO�����`�C(ڴr�YE�X�����jsK�T�~"Ȏ������Vv-=�__dG�2a]?jG̲Qm?j�c;՞�j�Q��b"��GmSl������[0�_eG������KMD�gt�.=��\���DT���-0��$V!C�9K�������<d �M9���l�T�Z�-�پx���	��ǌ��32�.����U�mױ��cU�zV�w�h���R+.7���q�<�1/F���;���RlH1W��TUR�%���JUf����s1�9J�����9��`�#J+�dh�^(mֹ�2���!5�r*���@�'a�A:��~ 5$
��c���1�v �1�h�� gt�`�h�XD5ց=�ɱ)Ȕ��U��4)��z�&～J���O) C.�,E"ͳ\<]O�]̞��X���ߖ_G)&K�L!c�J ��=3�`� �Ѡ	Sٝ�M4�hC��Hk`������L_O�N�I#����k�=KSnX���:W�p�I�D����ђp��n�6���qy��ղ�/
�I��x�w��;���'d��WW�	��R�;y���4��?���D�E&��x��x�(�A�x.!5�F��}��{�D��B��dL���S)�{y�l*�:��<��(���SԥX�h3�siȩ�ņ�j�˩%Q�t:)��l�PZ���ʚiJV�A��o���!��D:4jA��M˱�6P����DiN�V 9-�_h��v�I�Q@��H�m���������5ko$����h�^����KG��)Ӧ:� C�g`T�����r8m�rn!�or'�"}�aqgݙ�0`Bh�X�Gϲ��
@
��Q*�Ř�<;��
J$ �5k#�l�	N����J	4�h`�J���#���wvVE{l�2i����t��4��.�i�h��j�6���lwD,�h*�6�����y��R>h�P$��������KR��<�~C��tc�hCvu��QN	�}k)X��t�;��J<(����J5��ݳM^ ���[ѐ��R9~�=��]G ���`c��	R9VI��~mS=jK%�BKR9CE�����'|kl� mo�c����K��|�ܓ�Dp!����>ء>��䔠,�	*b��]�#�V�\HC:�|��opcG�iR����Yv5�eUBY�{(�B'G��/��՞6���R�0��~��N�q�RT�N�����A&�R�6�?���hv^O�hw}�1}��� 0"%��9�)@r��2�~�P]Ǳ�w���+
�|4w럀�`0R �H	����x��lZ��i��H��F���i~�PK
   ���X��/�   ί                  cirkitFile.jsonPK
   ���XWC��)�  � /             �   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   ���X� ���� 
� /             Q�  images/38cb4f51-bc72-4d24-b782-e5d855ce8001.pngPK
   ���X����+  J  /             �� images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   ���X��_8
  3
  /             � images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   ���X����H   C   /             �� images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   ���X��) oj /             *� images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
   �X�X#&g��x hz /             �
 images/a033a989-baef-4d73-a136-ed3ff270941b.pngPK
   ���X$7h�!  �!  /             �� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ���X~��a� ٮ /             � images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   ���X�'k�  �  /             �a images/e8452abc-1b33-4025-a556-b46ce3c60df1.pngPK
   �X�X1��	B6 �8 /             �x images/e9cc877d-5fca-438f-8a74-200c5bfeb6c1.pngPK
   ���XP��/�  ǽ  /             {� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ���X����G	  ~.               �a jsons/user_defined.jsonPK      �  Ik   